module fir2n (clk, rst, din[0], din[1], din[2], din[3], din[4], din[5], din[6], din[7], dout[0], dout[1], dout[2], dout[3], dout[4], dout[5], dout[6], dout[7]);

input clk;
input rst;
input din[0];
input din[1];
input din[2];
input din[3];
input din[4];
input din[5];
input din[6];
input din[7];
output dout[0];
output dout[1];
output dout[2];
output dout[3];
output dout[4];
output dout[5];
output dout[6];
output dout[7];

BUFX2 BUFX2_1 ( .A(clk2_clkout), .Y(clk2_clkout_hier0_bF_buf5) );
BUFX2 BUFX2_2 ( .A(clk2_clkout), .Y(clk2_clkout_hier0_bF_buf4) );
BUFX2 BUFX2_3 ( .A(clk2_clkout), .Y(clk2_clkout_hier0_bF_buf3) );
BUFX2 BUFX2_4 ( .A(clk2_clkout), .Y(clk2_clkout_hier0_bF_buf2) );
BUFX2 BUFX2_5 ( .A(clk2_clkout), .Y(clk2_clkout_hier0_bF_buf1) );
BUFX2 BUFX2_6 ( .A(clk2_clkout), .Y(clk2_clkout_hier0_bF_buf0) );
BUFX2 BUFX2_7 ( .A(counterup_counter_0_), .Y(counterup_counter_0_bF_buf3_) );
BUFX2 BUFX2_8 ( .A(counterup_counter_0_), .Y(counterup_counter_0_bF_buf2_) );
BUFX2 BUFX2_9 ( .A(counterup_counter_0_), .Y(counterup_counter_0_bF_buf1_) );
BUFX2 BUFX2_10 ( .A(counterup_counter_0_), .Y(counterup_counter_0_bF_buf0_) );
CLKBUF1 CLKBUF1_1 ( .A(clk2_clkout_hier0_bF_buf4), .Y(clk2_clkout_bF_buf41) );
CLKBUF1 CLKBUF1_2 ( .A(clk2_clkout_hier0_bF_buf1), .Y(clk2_clkout_bF_buf40) );
CLKBUF1 CLKBUF1_3 ( .A(clk2_clkout_hier0_bF_buf0), .Y(clk2_clkout_bF_buf39) );
CLKBUF1 CLKBUF1_4 ( .A(clk2_clkout_hier0_bF_buf5), .Y(clk2_clkout_bF_buf38) );
CLKBUF1 CLKBUF1_5 ( .A(clk2_clkout_hier0_bF_buf2), .Y(clk2_clkout_bF_buf37) );
CLKBUF1 CLKBUF1_6 ( .A(clk2_clkout_hier0_bF_buf1), .Y(clk2_clkout_bF_buf36) );
CLKBUF1 CLKBUF1_7 ( .A(clk2_clkout_hier0_bF_buf0), .Y(clk2_clkout_bF_buf35) );
CLKBUF1 CLKBUF1_8 ( .A(clk2_clkout_hier0_bF_buf2), .Y(clk2_clkout_bF_buf34) );
CLKBUF1 CLKBUF1_9 ( .A(clk2_clkout_hier0_bF_buf5), .Y(clk2_clkout_bF_buf33) );
CLKBUF1 CLKBUF1_10 ( .A(clk2_clkout_hier0_bF_buf1), .Y(clk2_clkout_bF_buf32) );
CLKBUF1 CLKBUF1_11 ( .A(clk2_clkout_hier0_bF_buf2), .Y(clk2_clkout_bF_buf31) );
CLKBUF1 CLKBUF1_12 ( .A(clk2_clkout_hier0_bF_buf1), .Y(clk2_clkout_bF_buf30) );
CLKBUF1 CLKBUF1_13 ( .A(clk2_clkout_hier0_bF_buf5), .Y(clk2_clkout_bF_buf29) );
CLKBUF1 CLKBUF1_14 ( .A(clk2_clkout_hier0_bF_buf1), .Y(clk2_clkout_bF_buf28) );
CLKBUF1 CLKBUF1_15 ( .A(clk2_clkout_hier0_bF_buf3), .Y(clk2_clkout_bF_buf27) );
CLKBUF1 CLKBUF1_16 ( .A(clk2_clkout_hier0_bF_buf4), .Y(clk2_clkout_bF_buf26) );
CLKBUF1 CLKBUF1_17 ( .A(clk2_clkout_hier0_bF_buf2), .Y(clk2_clkout_bF_buf25) );
CLKBUF1 CLKBUF1_18 ( .A(clk2_clkout_hier0_bF_buf3), .Y(clk2_clkout_bF_buf24) );
CLKBUF1 CLKBUF1_19 ( .A(clk2_clkout_hier0_bF_buf3), .Y(clk2_clkout_bF_buf23) );
CLKBUF1 CLKBUF1_20 ( .A(clk2_clkout_hier0_bF_buf1), .Y(clk2_clkout_bF_buf22) );
CLKBUF1 CLKBUF1_21 ( .A(clk2_clkout_hier0_bF_buf3), .Y(clk2_clkout_bF_buf21) );
CLKBUF1 CLKBUF1_22 ( .A(clk2_clkout_hier0_bF_buf0), .Y(clk2_clkout_bF_buf20) );
CLKBUF1 CLKBUF1_23 ( .A(clk2_clkout_hier0_bF_buf4), .Y(clk2_clkout_bF_buf19) );
CLKBUF1 CLKBUF1_24 ( .A(clk2_clkout_hier0_bF_buf4), .Y(clk2_clkout_bF_buf18) );
CLKBUF1 CLKBUF1_25 ( .A(clk2_clkout_hier0_bF_buf3), .Y(clk2_clkout_bF_buf17) );
CLKBUF1 CLKBUF1_26 ( .A(clk2_clkout_hier0_bF_buf2), .Y(clk2_clkout_bF_buf16) );
CLKBUF1 CLKBUF1_27 ( .A(clk2_clkout_hier0_bF_buf0), .Y(clk2_clkout_bF_buf15) );
CLKBUF1 CLKBUF1_28 ( .A(clk2_clkout_hier0_bF_buf5), .Y(clk2_clkout_bF_buf14) );
CLKBUF1 CLKBUF1_29 ( .A(clk2_clkout_hier0_bF_buf0), .Y(clk2_clkout_bF_buf13) );
CLKBUF1 CLKBUF1_30 ( .A(clk2_clkout_hier0_bF_buf4), .Y(clk2_clkout_bF_buf12) );
CLKBUF1 CLKBUF1_31 ( .A(clk2_clkout_hier0_bF_buf3), .Y(clk2_clkout_bF_buf11) );
CLKBUF1 CLKBUF1_32 ( .A(clk2_clkout_hier0_bF_buf3), .Y(clk2_clkout_bF_buf10) );
CLKBUF1 CLKBUF1_33 ( .A(clk2_clkout_hier0_bF_buf2), .Y(clk2_clkout_bF_buf9) );
CLKBUF1 CLKBUF1_34 ( .A(clk2_clkout_hier0_bF_buf1), .Y(clk2_clkout_bF_buf8) );
CLKBUF1 CLKBUF1_35 ( .A(clk2_clkout_hier0_bF_buf4), .Y(clk2_clkout_bF_buf7) );
CLKBUF1 CLKBUF1_36 ( .A(clk2_clkout_hier0_bF_buf2), .Y(clk2_clkout_bF_buf6) );
CLKBUF1 CLKBUF1_37 ( .A(clk2_clkout_hier0_bF_buf5), .Y(clk2_clkout_bF_buf5) );
CLKBUF1 CLKBUF1_38 ( .A(clk2_clkout_hier0_bF_buf5), .Y(clk2_clkout_bF_buf4) );
CLKBUF1 CLKBUF1_39 ( .A(clk2_clkout_hier0_bF_buf0), .Y(clk2_clkout_bF_buf3) );
CLKBUF1 CLKBUF1_40 ( .A(clk2_clkout_hier0_bF_buf0), .Y(clk2_clkout_bF_buf2) );
CLKBUF1 CLKBUF1_41 ( .A(clk2_clkout_hier0_bF_buf5), .Y(clk2_clkout_bF_buf1) );
CLKBUF1 CLKBUF1_42 ( .A(clk2_clkout_hier0_bF_buf4), .Y(clk2_clkout_bF_buf0) );
BUFX2 BUFX2_11 ( .A(_4_), .Y(_4__bF_buf3) );
BUFX2 BUFX2_12 ( .A(_4_), .Y(_4__bF_buf2) );
BUFX2 BUFX2_13 ( .A(_4_), .Y(_4__bF_buf1) );
BUFX2 BUFX2_14 ( .A(_4_), .Y(_4__bF_buf0) );
CLKBUF1 CLKBUF1_43 ( .A(clk), .Y(clk_bF_buf6) );
CLKBUF1 CLKBUF1_44 ( .A(clk), .Y(clk_bF_buf5) );
CLKBUF1 CLKBUF1_45 ( .A(clk), .Y(clk_bF_buf4) );
CLKBUF1 CLKBUF1_46 ( .A(clk), .Y(clk_bF_buf3) );
CLKBUF1 CLKBUF1_47 ( .A(clk), .Y(clk_bF_buf2) );
CLKBUF1 CLKBUF1_48 ( .A(clk), .Y(clk_bF_buf1) );
CLKBUF1 CLKBUF1_49 ( .A(clk), .Y(clk_bF_buf0) );
BUFX2 BUFX2_15 ( .A(_36_), .Y(_36__bF_buf3) );
BUFX2 BUFX2_16 ( .A(_36_), .Y(_36__bF_buf2) );
BUFX2 BUFX2_17 ( .A(_36_), .Y(_36__bF_buf1) );
BUFX2 BUFX2_18 ( .A(_36_), .Y(_36__bF_buf0) );
BUFX2 BUFX2_19 ( .A(_33_), .Y(_33__bF_buf3) );
BUFX2 BUFX2_20 ( .A(_33_), .Y(_33__bF_buf2) );
BUFX2 BUFX2_21 ( .A(_33_), .Y(_33__bF_buf1) );
BUFX2 BUFX2_22 ( .A(_33_), .Y(_33__bF_buf0) );
BUFX2 BUFX2_23 ( .A(_229_), .Y(_229__bF_buf3) );
BUFX2 BUFX2_24 ( .A(_229_), .Y(_229__bF_buf2) );
BUFX2 BUFX2_25 ( .A(_229_), .Y(_229__bF_buf1) );
BUFX2 BUFX2_26 ( .A(_229_), .Y(_229__bF_buf0) );
BUFX2 BUFX2_27 ( .A(_261_), .Y(_261__bF_buf3) );
BUFX2 BUFX2_28 ( .A(_261_), .Y(_261__bF_buf2) );
BUFX2 BUFX2_29 ( .A(_261_), .Y(_261__bF_buf1) );
BUFX2 BUFX2_30 ( .A(_261_), .Y(_261__bF_buf0) );
BUFX2 BUFX2_31 ( .A(_258_), .Y(_258__bF_buf3) );
BUFX2 BUFX2_32 ( .A(_258_), .Y(_258__bF_buf2) );
BUFX2 BUFX2_33 ( .A(_258_), .Y(_258__bF_buf1) );
BUFX2 BUFX2_34 ( .A(_258_), .Y(_258__bF_buf0) );
BUFX2 BUFX2_35 ( .A(rst), .Y(rst_bF_buf5) );
BUFX2 BUFX2_36 ( .A(rst), .Y(rst_bF_buf4) );
BUFX2 BUFX2_37 ( .A(rst), .Y(rst_bF_buf3) );
BUFX2 BUFX2_38 ( .A(rst), .Y(rst_bF_buf2) );
BUFX2 BUFX2_39 ( .A(rst), .Y(rst_bF_buf1) );
BUFX2 BUFX2_40 ( .A(rst), .Y(rst_bF_buf0) );
BUFX2 BUFX2_41 ( .A(_0_), .Y(_0__bF_buf10) );
BUFX2 BUFX2_42 ( .A(_0_), .Y(_0__bF_buf9) );
BUFX2 BUFX2_43 ( .A(_0_), .Y(_0__bF_buf8) );
BUFX2 BUFX2_44 ( .A(_0_), .Y(_0__bF_buf7) );
BUFX2 BUFX2_45 ( .A(_0_), .Y(_0__bF_buf6) );
BUFX2 BUFX2_46 ( .A(_0_), .Y(_0__bF_buf5) );
BUFX2 BUFX2_47 ( .A(_0_), .Y(_0__bF_buf4) );
BUFX2 BUFX2_48 ( .A(_0_), .Y(_0__bF_buf3) );
BUFX2 BUFX2_49 ( .A(_0_), .Y(_0__bF_buf2) );
BUFX2 BUFX2_50 ( .A(_0_), .Y(_0__bF_buf1) );
BUFX2 BUFX2_51 ( .A(_0_), .Y(_0__bF_buf0) );
BUFX2 BUFX2_52 ( .A(mac1_reset), .Y(mac1_reset_bF_buf3) );
BUFX2 BUFX2_53 ( .A(mac1_reset), .Y(mac1_reset_bF_buf2) );
BUFX2 BUFX2_54 ( .A(mac1_reset), .Y(mac1_reset_bF_buf1) );
BUFX2 BUFX2_55 ( .A(mac1_reset), .Y(mac1_reset_bF_buf0) );
BUFX2 BUFX2_56 ( .A(rom1_data_0_), .Y(rom1_data_0_bF_buf3_) );
BUFX2 BUFX2_57 ( .A(rom1_data_0_), .Y(rom1_data_0_bF_buf2_) );
BUFX2 BUFX2_58 ( .A(rom1_data_0_), .Y(rom1_data_0_bF_buf1_) );
BUFX2 BUFX2_59 ( .A(rom1_data_0_), .Y(rom1_data_0_bF_buf0_) );
BUFX2 BUFX2_60 ( .A(_225_), .Y(_225__bF_buf10) );
BUFX2 BUFX2_61 ( .A(_225_), .Y(_225__bF_buf9) );
BUFX2 BUFX2_62 ( .A(_225_), .Y(_225__bF_buf8) );
BUFX2 BUFX2_63 ( .A(_225_), .Y(_225__bF_buf7) );
BUFX2 BUFX2_64 ( .A(_225_), .Y(_225__bF_buf6) );
BUFX2 BUFX2_65 ( .A(_225_), .Y(_225__bF_buf5) );
BUFX2 BUFX2_66 ( .A(_225_), .Y(_225__bF_buf4) );
BUFX2 BUFX2_67 ( .A(_225_), .Y(_225__bF_buf3) );
BUFX2 BUFX2_68 ( .A(_225_), .Y(_225__bF_buf2) );
BUFX2 BUFX2_69 ( .A(_225_), .Y(_225__bF_buf1) );
BUFX2 BUFX2_70 ( .A(_225_), .Y(_225__bF_buf0) );
BUFX2 BUFX2_71 ( .A(reg3_dataout_0_), .Y(dout[0]) );
BUFX2 BUFX2_72 ( .A(reg3_dataout_1_), .Y(dout[1]) );
BUFX2 BUFX2_73 ( .A(reg3_dataout_2_), .Y(dout[2]) );
BUFX2 BUFX2_74 ( .A(reg3_dataout_3_), .Y(dout[3]) );
BUFX2 BUFX2_75 ( .A(reg3_dataout_4_), .Y(dout[4]) );
BUFX2 BUFX2_76 ( .A(reg3_dataout_5_), .Y(dout[5]) );
BUFX2 BUFX2_77 ( .A(reg3_dataout_6_), .Y(dout[6]) );
BUFX2 BUFX2_78 ( .A(reg3_dataout_7_), .Y(dout[7]) );
INVX1 INVX1_1 ( .A(asr1_rom_6__0_), .Y(_1_) );
INVX1 INVX1_2 ( .A(asr1_rom_5__0_), .Y(_2_) );
INVX1 INVX1_3 ( .A(counterup_counter_3_), .Y(_3_) );
AND2X2 AND2X2_1 ( .A(_3_), .B(counterup_counter_2_), .Y(_4_) );
INVX1 INVX1_4 ( .A(counterup_counter_1_), .Y(_5_) );
AND2X2 AND2X2_2 ( .A(_5_), .B(counterup_counter_0_bF_buf3_), .Y(_6_) );
NAND2X1 NAND2X1_1 ( .A(_4__bF_buf2), .B(_6_), .Y(_7_) );
NOR2X1 NOR2X1_1 ( .A(counterup_counter_0_bF_buf2_), .B(_5_), .Y(_8_) );
NAND2X1 NAND2X1_2 ( .A(_8_), .B(_4__bF_buf3), .Y(_9_) );
OAI22X1 OAI22X1_1 ( .A(_1_), .B(_9_), .C(_2_), .D(_7_), .Y(_10_) );
INVX1 INVX1_5 ( .A(asr1_rom_10__0_), .Y(_11_) );
INVX1 INVX1_6 ( .A(asr1_rom_9__0_), .Y(_12_) );
NOR2X1 NOR2X1_2 ( .A(counterup_counter_2_), .B(_3_), .Y(_13_) );
NAND2X1 NAND2X1_3 ( .A(_13_), .B(_6_), .Y(_14_) );
NAND2X1 NAND2X1_4 ( .A(_8_), .B(_13_), .Y(_15_) );
OAI22X1 OAI22X1_2 ( .A(_11_), .B(_15_), .C(_12_), .D(_14_), .Y(_16_) );
NOR2X1 NOR2X1_3 ( .A(_16_), .B(_10_), .Y(_17_) );
INVX1 INVX1_7 ( .A(asr1_rom_2__0_), .Y(_18_) );
INVX1 INVX1_8 ( .A(asr1_rom_1__0_), .Y(_19_) );
NOR2X1 NOR2X1_4 ( .A(counterup_counter_3_), .B(counterup_counter_2_), .Y(_20_) );
NAND2X1 NAND2X1_5 ( .A(_20_), .B(_6_), .Y(_21_) );
NAND2X1 NAND2X1_6 ( .A(_20_), .B(_8_), .Y(_22_) );
OAI22X1 OAI22X1_3 ( .A(_18_), .B(_22_), .C(_19_), .D(_21_), .Y(_23_) );
INVX1 INVX1_9 ( .A(asr1_rom_14__0_), .Y(_24_) );
NAND2X1 NAND2X1_7 ( .A(counterup_counter_0_bF_buf1_), .B(_5_), .Y(_25_) );
NAND2X1 NAND2X1_8 ( .A(counterup_counter_3_), .B(counterup_counter_2_), .Y(_26_) );
NOR2X1 NOR2X1_5 ( .A(_26_), .B(_25_), .Y(_27_) );
NAND2X1 NAND2X1_9 ( .A(asr1_rom_13__0_), .B(_27_), .Y(_28_) );
AND2X2 AND2X2_3 ( .A(counterup_counter_3_), .B(counterup_counter_2_), .Y(_29_) );
NAND2X1 NAND2X1_10 ( .A(_29_), .B(_8_), .Y(_30_) );
OAI21X1 OAI21X1_1 ( .A(_24_), .B(_30_), .C(_28_), .Y(_31_) );
NOR2X1 NOR2X1_6 ( .A(_23_), .B(_31_), .Y(_32_) );
AND2X2 AND2X2_4 ( .A(counterup_counter_1_), .B(counterup_counter_0_bF_buf0_), .Y(_33_) );
AND2X2 AND2X2_5 ( .A(_33__bF_buf3), .B(_20_), .Y(_34_) );
NAND2X1 NAND2X1_11 ( .A(asr1_rom_3__0_), .B(_34_), .Y(_35_) );
NOR2X1 NOR2X1_7 ( .A(counterup_counter_1_), .B(counterup_counter_0_bF_buf3_), .Y(_36_) );
NAND3X1 NAND3X1_1 ( .A(asr1_rom_4__0_), .B(_36__bF_buf2), .C(_4__bF_buf0), .Y(_37_) );
NAND3X1 NAND3X1_2 ( .A(asr1_rom_0__0_), .B(_20_), .C(_36__bF_buf2), .Y(_38_) );
NAND3X1 NAND3X1_3 ( .A(asr1_en_0_), .B(_29_), .C(_33__bF_buf2), .Y(_39_) );
AND2X2 AND2X2_6 ( .A(_39_), .B(_38_), .Y(_40_) );
NAND3X1 NAND3X1_4 ( .A(_35_), .B(_37_), .C(_40_), .Y(_41_) );
NAND3X1 NAND3X1_5 ( .A(asr1_rom_7__0_), .B(_33__bF_buf0), .C(_4__bF_buf3), .Y(_42_) );
NAND3X1 NAND3X1_6 ( .A(asr1_rom_8__0_), .B(_36__bF_buf2), .C(_13_), .Y(_43_) );
NAND2X1 NAND2X1_12 ( .A(counterup_counter_1_), .B(counterup_counter_0_bF_buf2_), .Y(_44_) );
NOR3X1 NOR3X1_1 ( .A(counterup_counter_2_), .B(_3_), .C(_44_), .Y(_45_) );
NOR3X1 NOR3X1_2 ( .A(counterup_counter_1_), .B(counterup_counter_0_bF_buf1_), .C(_26_), .Y(_46_) );
AOI22X1 AOI22X1_1 ( .A(_46_), .B(asr1_rom_12__0_), .C(asr1_rom_11__0_), .D(_45_), .Y(_47_) );
NAND3X1 NAND3X1_7 ( .A(_42_), .B(_43_), .C(_47_), .Y(_48_) );
NOR2X1 NOR2X1_8 ( .A(_41_), .B(_48_), .Y(_49_) );
NAND3X1 NAND3X1_8 ( .A(_17_), .B(_32_), .C(_49_), .Y(asr1_dataout_0_) );
INVX1 INVX1_10 ( .A(asr1_rom_6__1_), .Y(_50_) );
INVX1 INVX1_11 ( .A(asr1_rom_5__1_), .Y(_51_) );
OAI22X1 OAI22X1_4 ( .A(_50_), .B(_9_), .C(_51_), .D(_7_), .Y(_52_) );
INVX1 INVX1_12 ( .A(asr1_rom_10__1_), .Y(_53_) );
INVX1 INVX1_13 ( .A(asr1_rom_9__1_), .Y(_54_) );
OAI22X1 OAI22X1_5 ( .A(_53_), .B(_15_), .C(_54_), .D(_14_), .Y(_55_) );
NOR2X1 NOR2X1_9 ( .A(_55_), .B(_52_), .Y(_56_) );
INVX1 INVX1_14 ( .A(asr1_rom_2__1_), .Y(_57_) );
INVX1 INVX1_15 ( .A(asr1_rom_1__1_), .Y(_58_) );
OAI22X1 OAI22X1_6 ( .A(_57_), .B(_22_), .C(_58_), .D(_21_), .Y(_59_) );
INVX1 INVX1_16 ( .A(asr1_rom_14__1_), .Y(_60_) );
NAND2X1 NAND2X1_13 ( .A(asr1_rom_13__1_), .B(_27_), .Y(_61_) );
OAI21X1 OAI21X1_2 ( .A(_60_), .B(_30_), .C(_61_), .Y(_62_) );
NOR2X1 NOR2X1_10 ( .A(_59_), .B(_62_), .Y(_63_) );
NAND2X1 NAND2X1_14 ( .A(asr1_rom_3__1_), .B(_34_), .Y(_64_) );
NAND3X1 NAND3X1_9 ( .A(asr1_rom_4__1_), .B(_36__bF_buf1), .C(_4__bF_buf2), .Y(_65_) );
NAND3X1 NAND3X1_10 ( .A(asr1_rom_0__1_), .B(_20_), .C(_36__bF_buf0), .Y(_66_) );
NAND3X1 NAND3X1_11 ( .A(asr1_en_1_), .B(_29_), .C(_33__bF_buf1), .Y(_67_) );
AND2X2 AND2X2_7 ( .A(_67_), .B(_66_), .Y(_68_) );
NAND3X1 NAND3X1_12 ( .A(_64_), .B(_65_), .C(_68_), .Y(_69_) );
NAND3X1 NAND3X1_13 ( .A(asr1_rom_7__1_), .B(_33__bF_buf3), .C(_4__bF_buf1), .Y(_70_) );
NAND3X1 NAND3X1_14 ( .A(asr1_rom_8__1_), .B(_36__bF_buf3), .C(_13_), .Y(_71_) );
AOI22X1 AOI22X1_2 ( .A(_46_), .B(asr1_rom_12__1_), .C(asr1_rom_11__1_), .D(_45_), .Y(_72_) );
NAND3X1 NAND3X1_15 ( .A(_70_), .B(_71_), .C(_72_), .Y(_73_) );
NOR2X1 NOR2X1_11 ( .A(_69_), .B(_73_), .Y(_74_) );
NAND3X1 NAND3X1_16 ( .A(_56_), .B(_63_), .C(_74_), .Y(asr1_dataout_1_) );
INVX1 INVX1_17 ( .A(asr1_rom_6__2_), .Y(_75_) );
INVX1 INVX1_18 ( .A(asr1_rom_5__2_), .Y(_76_) );
OAI22X1 OAI22X1_7 ( .A(_75_), .B(_9_), .C(_76_), .D(_7_), .Y(_77_) );
INVX1 INVX1_19 ( .A(asr1_rom_10__2_), .Y(_78_) );
INVX1 INVX1_20 ( .A(asr1_rom_9__2_), .Y(_79_) );
OAI22X1 OAI22X1_8 ( .A(_78_), .B(_15_), .C(_79_), .D(_14_), .Y(_80_) );
NOR2X1 NOR2X1_12 ( .A(_80_), .B(_77_), .Y(_81_) );
INVX1 INVX1_21 ( .A(asr1_rom_2__2_), .Y(_82_) );
INVX1 INVX1_22 ( .A(asr1_rom_1__2_), .Y(_83_) );
OAI22X1 OAI22X1_9 ( .A(_82_), .B(_22_), .C(_83_), .D(_21_), .Y(_84_) );
INVX1 INVX1_23 ( .A(asr1_rom_14__2_), .Y(_85_) );
NAND2X1 NAND2X1_15 ( .A(asr1_rom_13__2_), .B(_27_), .Y(_86_) );
OAI21X1 OAI21X1_3 ( .A(_85_), .B(_30_), .C(_86_), .Y(_87_) );
NOR2X1 NOR2X1_13 ( .A(_84_), .B(_87_), .Y(_88_) );
NAND2X1 NAND2X1_16 ( .A(asr1_rom_3__2_), .B(_34_), .Y(_89_) );
NAND3X1 NAND3X1_17 ( .A(asr1_rom_4__2_), .B(_36__bF_buf2), .C(_4__bF_buf3), .Y(_90_) );
NAND3X1 NAND3X1_18 ( .A(asr1_rom_0__2_), .B(_20_), .C(_36__bF_buf2), .Y(_91_) );
NAND3X1 NAND3X1_19 ( .A(asr1_en_2_), .B(_29_), .C(_33__bF_buf2), .Y(_92_) );
AND2X2 AND2X2_8 ( .A(_92_), .B(_91_), .Y(_93_) );
NAND3X1 NAND3X1_20 ( .A(_89_), .B(_90_), .C(_93_), .Y(_94_) );
NAND3X1 NAND3X1_21 ( .A(asr1_rom_7__2_), .B(_33__bF_buf0), .C(_4__bF_buf3), .Y(_95_) );
NAND3X1 NAND3X1_22 ( .A(asr1_rom_8__2_), .B(_36__bF_buf0), .C(_13_), .Y(_96_) );
AOI22X1 AOI22X1_3 ( .A(_46_), .B(asr1_rom_12__2_), .C(asr1_rom_11__2_), .D(_45_), .Y(_97_) );
NAND3X1 NAND3X1_23 ( .A(_95_), .B(_96_), .C(_97_), .Y(_98_) );
NOR2X1 NOR2X1_14 ( .A(_94_), .B(_98_), .Y(_99_) );
NAND3X1 NAND3X1_24 ( .A(_81_), .B(_88_), .C(_99_), .Y(asr1_dataout_2_) );
INVX1 INVX1_24 ( .A(asr1_rom_6__3_), .Y(_100_) );
INVX1 INVX1_25 ( .A(asr1_rom_5__3_), .Y(_101_) );
OAI22X1 OAI22X1_10 ( .A(_100_), .B(_9_), .C(_101_), .D(_7_), .Y(_102_) );
INVX1 INVX1_26 ( .A(asr1_rom_10__3_), .Y(_103_) );
INVX1 INVX1_27 ( .A(asr1_rom_9__3_), .Y(_104_) );
OAI22X1 OAI22X1_11 ( .A(_103_), .B(_15_), .C(_104_), .D(_14_), .Y(_105_) );
NOR2X1 NOR2X1_15 ( .A(_105_), .B(_102_), .Y(_106_) );
INVX1 INVX1_28 ( .A(asr1_rom_2__3_), .Y(_107_) );
INVX1 INVX1_29 ( .A(asr1_rom_1__3_), .Y(_108_) );
OAI22X1 OAI22X1_12 ( .A(_107_), .B(_22_), .C(_108_), .D(_21_), .Y(_109_) );
INVX1 INVX1_30 ( .A(asr1_rom_14__3_), .Y(_110_) );
NAND2X1 NAND2X1_17 ( .A(asr1_rom_13__3_), .B(_27_), .Y(_111_) );
OAI21X1 OAI21X1_4 ( .A(_110_), .B(_30_), .C(_111_), .Y(_112_) );
NOR2X1 NOR2X1_16 ( .A(_109_), .B(_112_), .Y(_113_) );
NAND2X1 NAND2X1_18 ( .A(asr1_rom_3__3_), .B(_34_), .Y(_114_) );
NAND3X1 NAND3X1_25 ( .A(asr1_rom_4__3_), .B(_36__bF_buf1), .C(_4__bF_buf2), .Y(_115_) );
NAND3X1 NAND3X1_26 ( .A(asr1_rom_0__3_), .B(_20_), .C(_36__bF_buf1), .Y(_116_) );
NAND3X1 NAND3X1_27 ( .A(asr1_en_3_), .B(_29_), .C(_33__bF_buf1), .Y(_117_) );
AND2X2 AND2X2_9 ( .A(_117_), .B(_116_), .Y(_118_) );
NAND3X1 NAND3X1_28 ( .A(_114_), .B(_115_), .C(_118_), .Y(_119_) );
NAND3X1 NAND3X1_29 ( .A(asr1_rom_7__3_), .B(_33__bF_buf1), .C(_4__bF_buf2), .Y(_120_) );
NAND3X1 NAND3X1_30 ( .A(asr1_rom_8__3_), .B(_36__bF_buf0), .C(_13_), .Y(_121_) );
AOI22X1 AOI22X1_4 ( .A(_46_), .B(asr1_rom_12__3_), .C(asr1_rom_11__3_), .D(_45_), .Y(_122_) );
NAND3X1 NAND3X1_31 ( .A(_120_), .B(_121_), .C(_122_), .Y(_123_) );
NOR2X1 NOR2X1_17 ( .A(_119_), .B(_123_), .Y(_124_) );
NAND3X1 NAND3X1_32 ( .A(_106_), .B(_113_), .C(_124_), .Y(asr1_dataout_3_) );
INVX1 INVX1_31 ( .A(asr1_rom_6__4_), .Y(_125_) );
INVX1 INVX1_32 ( .A(asr1_rom_5__4_), .Y(_126_) );
OAI22X1 OAI22X1_13 ( .A(_125_), .B(_9_), .C(_126_), .D(_7_), .Y(_127_) );
INVX1 INVX1_33 ( .A(asr1_rom_10__4_), .Y(_128_) );
INVX1 INVX1_34 ( .A(asr1_rom_9__4_), .Y(_129_) );
OAI22X1 OAI22X1_14 ( .A(_128_), .B(_15_), .C(_129_), .D(_14_), .Y(_130_) );
NOR2X1 NOR2X1_18 ( .A(_130_), .B(_127_), .Y(_131_) );
INVX1 INVX1_35 ( .A(asr1_rom_2__4_), .Y(_132_) );
INVX1 INVX1_36 ( .A(asr1_rom_1__4_), .Y(_133_) );
OAI22X1 OAI22X1_15 ( .A(_132_), .B(_22_), .C(_133_), .D(_21_), .Y(_134_) );
INVX1 INVX1_37 ( .A(asr1_rom_14__4_), .Y(_135_) );
NAND2X1 NAND2X1_19 ( .A(asr1_rom_13__4_), .B(_27_), .Y(_136_) );
OAI21X1 OAI21X1_5 ( .A(_135_), .B(_30_), .C(_136_), .Y(_137_) );
NOR2X1 NOR2X1_19 ( .A(_134_), .B(_137_), .Y(_138_) );
NAND2X1 NAND2X1_20 ( .A(asr1_rom_3__4_), .B(_34_), .Y(_139_) );
NAND3X1 NAND3X1_33 ( .A(asr1_rom_4__4_), .B(_36__bF_buf3), .C(_4__bF_buf0), .Y(_140_) );
NAND3X1 NAND3X1_34 ( .A(asr1_rom_0__4_), .B(_20_), .C(_36__bF_buf3), .Y(_141_) );
NAND3X1 NAND3X1_35 ( .A(asr1_en_4_), .B(_29_), .C(_33__bF_buf2), .Y(_142_) );
AND2X2 AND2X2_10 ( .A(_142_), .B(_141_), .Y(_143_) );
NAND3X1 NAND3X1_36 ( .A(_139_), .B(_140_), .C(_143_), .Y(_144_) );
NAND3X1 NAND3X1_37 ( .A(asr1_rom_7__4_), .B(_33__bF_buf2), .C(_4__bF_buf0), .Y(_145_) );
NAND3X1 NAND3X1_38 ( .A(asr1_rom_8__4_), .B(_36__bF_buf2), .C(_13_), .Y(_146_) );
AOI22X1 AOI22X1_5 ( .A(_46_), .B(asr1_rom_12__4_), .C(asr1_rom_11__4_), .D(_45_), .Y(_147_) );
NAND3X1 NAND3X1_39 ( .A(_145_), .B(_146_), .C(_147_), .Y(_148_) );
NOR2X1 NOR2X1_20 ( .A(_144_), .B(_148_), .Y(_149_) );
NAND3X1 NAND3X1_40 ( .A(_131_), .B(_138_), .C(_149_), .Y(asr1_dataout_4_) );
INVX1 INVX1_38 ( .A(asr1_rom_6__5_), .Y(_150_) );
INVX1 INVX1_39 ( .A(asr1_rom_5__5_), .Y(_151_) );
OAI22X1 OAI22X1_16 ( .A(_150_), .B(_9_), .C(_151_), .D(_7_), .Y(_152_) );
INVX1 INVX1_40 ( .A(asr1_rom_10__5_), .Y(_153_) );
INVX1 INVX1_41 ( .A(asr1_rom_9__5_), .Y(_154_) );
OAI22X1 OAI22X1_17 ( .A(_153_), .B(_15_), .C(_154_), .D(_14_), .Y(_155_) );
NOR2X1 NOR2X1_21 ( .A(_155_), .B(_152_), .Y(_156_) );
INVX1 INVX1_42 ( .A(asr1_rom_2__5_), .Y(_157_) );
INVX1 INVX1_43 ( .A(asr1_rom_1__5_), .Y(_158_) );
OAI22X1 OAI22X1_18 ( .A(_157_), .B(_22_), .C(_158_), .D(_21_), .Y(_159_) );
INVX1 INVX1_44 ( .A(asr1_rom_14__5_), .Y(_160_) );
NAND2X1 NAND2X1_21 ( .A(asr1_rom_13__5_), .B(_27_), .Y(_161_) );
OAI21X1 OAI21X1_6 ( .A(_160_), .B(_30_), .C(_161_), .Y(_162_) );
NOR2X1 NOR2X1_22 ( .A(_159_), .B(_162_), .Y(_163_) );
NAND2X1 NAND2X1_22 ( .A(asr1_rom_3__5_), .B(_34_), .Y(_164_) );
NAND3X1 NAND3X1_41 ( .A(asr1_rom_4__5_), .B(_36__bF_buf0), .C(_4__bF_buf3), .Y(_165_) );
NAND3X1 NAND3X1_42 ( .A(asr1_rom_0__5_), .B(_20_), .C(_36__bF_buf0), .Y(_166_) );
NAND3X1 NAND3X1_43 ( .A(asr1_en_5_), .B(_29_), .C(_33__bF_buf0), .Y(_167_) );
AND2X2 AND2X2_11 ( .A(_167_), .B(_166_), .Y(_168_) );
NAND3X1 NAND3X1_44 ( .A(_164_), .B(_165_), .C(_168_), .Y(_169_) );
NAND3X1 NAND3X1_45 ( .A(asr1_rom_7__5_), .B(_33__bF_buf3), .C(_4__bF_buf1), .Y(_170_) );
NAND3X1 NAND3X1_46 ( .A(asr1_rom_8__5_), .B(_36__bF_buf3), .C(_13_), .Y(_171_) );
AOI22X1 AOI22X1_6 ( .A(_46_), .B(asr1_rom_12__5_), .C(asr1_rom_11__5_), .D(_45_), .Y(_172_) );
NAND3X1 NAND3X1_47 ( .A(_170_), .B(_171_), .C(_172_), .Y(_173_) );
NOR2X1 NOR2X1_23 ( .A(_169_), .B(_173_), .Y(_174_) );
NAND3X1 NAND3X1_48 ( .A(_156_), .B(_163_), .C(_174_), .Y(asr1_dataout_5_) );
INVX1 INVX1_45 ( .A(asr1_rom_6__6_), .Y(_175_) );
INVX1 INVX1_46 ( .A(asr1_rom_5__6_), .Y(_176_) );
OAI22X1 OAI22X1_19 ( .A(_175_), .B(_9_), .C(_176_), .D(_7_), .Y(_177_) );
INVX1 INVX1_47 ( .A(asr1_rom_10__6_), .Y(_178_) );
INVX1 INVX1_48 ( .A(asr1_rom_9__6_), .Y(_179_) );
OAI22X1 OAI22X1_20 ( .A(_178_), .B(_15_), .C(_179_), .D(_14_), .Y(_180_) );
NOR2X1 NOR2X1_24 ( .A(_180_), .B(_177_), .Y(_181_) );
INVX1 INVX1_49 ( .A(asr1_rom_2__6_), .Y(_182_) );
INVX1 INVX1_50 ( .A(asr1_rom_1__6_), .Y(_183_) );
OAI22X1 OAI22X1_21 ( .A(_182_), .B(_22_), .C(_183_), .D(_21_), .Y(_184_) );
INVX1 INVX1_51 ( .A(asr1_rom_14__6_), .Y(_185_) );
NAND2X1 NAND2X1_23 ( .A(asr1_rom_13__6_), .B(_27_), .Y(_186_) );
OAI21X1 OAI21X1_7 ( .A(_185_), .B(_30_), .C(_186_), .Y(_187_) );
NOR2X1 NOR2X1_25 ( .A(_184_), .B(_187_), .Y(_188_) );
NAND2X1 NAND2X1_24 ( .A(asr1_rom_3__6_), .B(_34_), .Y(_189_) );
NAND3X1 NAND3X1_49 ( .A(asr1_rom_4__6_), .B(_36__bF_buf1), .C(_4__bF_buf1), .Y(_190_) );
NAND3X1 NAND3X1_50 ( .A(asr1_rom_0__6_), .B(_20_), .C(_36__bF_buf0), .Y(_191_) );
NAND3X1 NAND3X1_51 ( .A(asr1_en_6_), .B(_29_), .C(_33__bF_buf0), .Y(_192_) );
AND2X2 AND2X2_12 ( .A(_192_), .B(_191_), .Y(_193_) );
NAND3X1 NAND3X1_52 ( .A(_189_), .B(_190_), .C(_193_), .Y(_194_) );
NAND3X1 NAND3X1_53 ( .A(asr1_rom_7__6_), .B(_33__bF_buf3), .C(_4__bF_buf1), .Y(_195_) );
NAND3X1 NAND3X1_54 ( .A(asr1_rom_8__6_), .B(_36__bF_buf3), .C(_13_), .Y(_196_) );
AOI22X1 AOI22X1_7 ( .A(_46_), .B(asr1_rom_12__6_), .C(asr1_rom_11__6_), .D(_45_), .Y(_197_) );
NAND3X1 NAND3X1_55 ( .A(_195_), .B(_196_), .C(_197_), .Y(_198_) );
NOR2X1 NOR2X1_26 ( .A(_194_), .B(_198_), .Y(_199_) );
NAND3X1 NAND3X1_56 ( .A(_181_), .B(_188_), .C(_199_), .Y(asr1_dataout_6_) );
INVX1 INVX1_52 ( .A(asr1_rom_6__7_), .Y(_200_) );
INVX1 INVX1_53 ( .A(asr1_rom_5__7_), .Y(_201_) );
OAI22X1 OAI22X1_22 ( .A(_200_), .B(_9_), .C(_201_), .D(_7_), .Y(_202_) );
INVX1 INVX1_54 ( .A(asr1_rom_10__7_), .Y(_203_) );
INVX1 INVX1_55 ( .A(asr1_rom_9__7_), .Y(_204_) );
OAI22X1 OAI22X1_23 ( .A(_203_), .B(_15_), .C(_204_), .D(_14_), .Y(_205_) );
NOR2X1 NOR2X1_27 ( .A(_205_), .B(_202_), .Y(_206_) );
INVX1 INVX1_56 ( .A(asr1_rom_2__7_), .Y(_207_) );
INVX1 INVX1_57 ( .A(asr1_rom_1__7_), .Y(_208_) );
OAI22X1 OAI22X1_24 ( .A(_207_), .B(_22_), .C(_208_), .D(_21_), .Y(_209_) );
INVX1 INVX1_58 ( .A(asr1_rom_14__7_), .Y(_210_) );
NAND2X1 NAND2X1_25 ( .A(asr1_rom_13__7_), .B(_27_), .Y(_211_) );
OAI21X1 OAI21X1_8 ( .A(_210_), .B(_30_), .C(_211_), .Y(_212_) );
NOR2X1 NOR2X1_28 ( .A(_209_), .B(_212_), .Y(_213_) );
NAND2X1 NAND2X1_26 ( .A(asr1_rom_3__7_), .B(_34_), .Y(_214_) );
NAND3X1 NAND3X1_57 ( .A(asr1_rom_4__7_), .B(_36__bF_buf1), .C(_4__bF_buf2), .Y(_215_) );
NAND3X1 NAND3X1_58 ( .A(asr1_rom_0__7_), .B(_20_), .C(_36__bF_buf1), .Y(_216_) );
NAND3X1 NAND3X1_59 ( .A(asr1_en_7_), .B(_29_), .C(_33__bF_buf1), .Y(_217_) );
AND2X2 AND2X2_13 ( .A(_217_), .B(_216_), .Y(_218_) );
NAND3X1 NAND3X1_60 ( .A(_214_), .B(_215_), .C(_218_), .Y(_219_) );
NAND3X1 NAND3X1_61 ( .A(asr1_rom_7__7_), .B(_33__bF_buf3), .C(_4__bF_buf0), .Y(_220_) );
NAND3X1 NAND3X1_62 ( .A(asr1_rom_8__7_), .B(_36__bF_buf3), .C(_13_), .Y(_221_) );
AOI22X1 AOI22X1_8 ( .A(_46_), .B(asr1_rom_12__7_), .C(asr1_rom_11__7_), .D(_45_), .Y(_222_) );
NAND3X1 NAND3X1_63 ( .A(_220_), .B(_221_), .C(_222_), .Y(_223_) );
NOR2X1 NOR2X1_29 ( .A(_219_), .B(_223_), .Y(_224_) );
NAND3X1 NAND3X1_64 ( .A(_206_), .B(_213_), .C(_224_), .Y(asr1_dataout_7_) );
INVX1 INVX1_59 ( .A(rst_bF_buf5), .Y(_0_) );
DFFSR DFFSR_1 ( .CLK(clk2_clkout_bF_buf23), .D(reg1_dataout_0_), .Q(asr1_rom_0__0_), .R(_0__bF_buf8), .S(1'b1) );
DFFSR DFFSR_2 ( .CLK(clk2_clkout_bF_buf14), .D(reg1_dataout_1_), .Q(asr1_rom_0__1_), .R(_0__bF_buf5), .S(1'b1) );
DFFSR DFFSR_3 ( .CLK(clk2_clkout_bF_buf41), .D(reg1_dataout_2_), .Q(asr1_rom_0__2_), .R(_0__bF_buf9), .S(1'b1) );
DFFSR DFFSR_4 ( .CLK(clk2_clkout_bF_buf38), .D(reg1_dataout_3_), .Q(asr1_rom_0__3_), .R(_0__bF_buf1), .S(1'b1) );
DFFSR DFFSR_5 ( .CLK(clk2_clkout_bF_buf12), .D(reg1_dataout_4_), .Q(asr1_rom_0__4_), .R(_0__bF_buf0), .S(1'b1) );
DFFSR DFFSR_6 ( .CLK(clk2_clkout_bF_buf14), .D(reg1_dataout_5_), .Q(asr1_rom_0__5_), .R(_0__bF_buf5), .S(1'b1) );
DFFSR DFFSR_7 ( .CLK(clk2_clkout_bF_buf33), .D(reg1_dataout_6_), .Q(asr1_rom_0__6_), .R(_0__bF_buf7), .S(1'b1) );
DFFSR DFFSR_8 ( .CLK(clk2_clkout_bF_buf29), .D(reg1_dataout_7_), .Q(asr1_rom_0__7_), .R(_0__bF_buf1), .S(1'b1) );
DFFSR DFFSR_9 ( .CLK(clk2_clkout_bF_buf16), .D(asr1_rom_6__0_), .Q(asr1_rom_7__0_), .R(_0__bF_buf4), .S(1'b1) );
DFFSR DFFSR_10 ( .CLK(clk2_clkout_bF_buf4), .D(asr1_rom_6__1_), .Q(asr1_rom_7__1_), .R(_0__bF_buf6), .S(1'b1) );
DFFSR DFFSR_11 ( .CLK(clk2_clkout_bF_buf34), .D(asr1_rom_6__2_), .Q(asr1_rom_7__2_), .R(_0__bF_buf8), .S(1'b1) );
DFFSR DFFSR_12 ( .CLK(clk2_clkout_bF_buf29), .D(asr1_rom_6__3_), .Q(asr1_rom_7__3_), .R(_0__bF_buf1), .S(1'b1) );
DFFSR DFFSR_13 ( .CLK(clk2_clkout_bF_buf16), .D(asr1_rom_6__4_), .Q(asr1_rom_7__4_), .R(_0__bF_buf3), .S(1'b1) );
DFFSR DFFSR_14 ( .CLK(clk2_clkout_bF_buf6), .D(asr1_rom_6__5_), .Q(asr1_rom_7__5_), .R(_0__bF_buf7), .S(1'b1) );
DFFSR DFFSR_15 ( .CLK(clk2_clkout_bF_buf5), .D(asr1_rom_6__6_), .Q(asr1_rom_7__6_), .R(_0__bF_buf6), .S(1'b1) );
DFFSR DFFSR_16 ( .CLK(clk2_clkout_bF_buf33), .D(asr1_rom_6__7_), .Q(asr1_rom_7__7_), .R(_0__bF_buf4), .S(1'b1) );
DFFSR DFFSR_17 ( .CLK(clk2_clkout_bF_buf35), .D(asr1_rom_1__0_), .Q(asr1_rom_2__0_), .R(_0__bF_buf9), .S(1'b1) );
DFFSR DFFSR_18 ( .CLK(clk2_clkout_bF_buf9), .D(asr1_rom_1__1_), .Q(asr1_rom_2__1_), .R(_0__bF_buf7), .S(1'b1) );
DFFSR DFFSR_19 ( .CLK(clk2_clkout_bF_buf35), .D(asr1_rom_1__2_), .Q(asr1_rom_2__2_), .R(_0__bF_buf9), .S(1'b1) );
DFFSR DFFSR_20 ( .CLK(clk2_clkout_bF_buf38), .D(asr1_rom_1__3_), .Q(asr1_rom_2__3_), .R(_0__bF_buf1), .S(1'b1) );
DFFSR DFFSR_21 ( .CLK(clk2_clkout_bF_buf7), .D(asr1_rom_1__4_), .Q(asr1_rom_2__4_), .R(_0__bF_buf0), .S(1'b1) );
DFFSR DFFSR_22 ( .CLK(clk2_clkout_bF_buf1), .D(asr1_rom_1__5_), .Q(asr1_rom_2__5_), .R(_0__bF_buf5), .S(1'b1) );
DFFSR DFFSR_23 ( .CLK(clk2_clkout_bF_buf24), .D(asr1_rom_1__6_), .Q(asr1_rom_2__6_), .R(_0__bF_buf8), .S(1'b1) );
DFFSR DFFSR_24 ( .CLK(clk2_clkout_bF_buf14), .D(asr1_rom_1__7_), .Q(asr1_rom_2__7_), .R(_0__bF_buf5), .S(1'b1) );
DFFSR DFFSR_25 ( .CLK(clk2_clkout_bF_buf35), .D(asr1_rom_0__0_), .Q(asr1_rom_1__0_), .R(_0__bF_buf9), .S(1'b1) );
DFFSR DFFSR_26 ( .CLK(clk2_clkout_bF_buf1), .D(asr1_rom_0__1_), .Q(asr1_rom_1__1_), .R(_0__bF_buf5), .S(1'b1) );
DFFSR DFFSR_27 ( .CLK(clk2_clkout_bF_buf41), .D(asr1_rom_0__2_), .Q(asr1_rom_1__2_), .R(_0__bF_buf9), .S(1'b1) );
DFFSR DFFSR_28 ( .CLK(clk2_clkout_bF_buf29), .D(asr1_rom_0__3_), .Q(asr1_rom_1__3_), .R(_0__bF_buf5), .S(1'b1) );
DFFSR DFFSR_29 ( .CLK(clk2_clkout_bF_buf18), .D(asr1_rom_0__4_), .Q(asr1_rom_1__4_), .R(_0__bF_buf0), .S(1'b1) );
DFFSR DFFSR_30 ( .CLK(clk2_clkout_bF_buf1), .D(asr1_rom_0__5_), .Q(asr1_rom_1__5_), .R(_0__bF_buf5), .S(1'b1) );
DFFSR DFFSR_31 ( .CLK(clk2_clkout_bF_buf33), .D(asr1_rom_0__6_), .Q(asr1_rom_1__6_), .R(_0__bF_buf4), .S(1'b1) );
DFFSR DFFSR_32 ( .CLK(clk2_clkout_bF_buf29), .D(asr1_rom_0__7_), .Q(asr1_rom_1__7_), .R(_0__bF_buf5), .S(1'b1) );
DFFSR DFFSR_33 ( .CLK(clk2_clkout_bF_buf35), .D(asr1_rom_2__0_), .Q(asr1_rom_3__0_), .R(_0__bF_buf9), .S(1'b1) );
DFFSR DFFSR_34 ( .CLK(clk2_clkout_bF_buf10), .D(asr1_rom_2__1_), .Q(asr1_rom_3__1_), .R(_0__bF_buf8), .S(1'b1) );
DFFSR DFFSR_35 ( .CLK(clk2_clkout_bF_buf26), .D(asr1_rom_2__2_), .Q(asr1_rom_3__2_), .R(_0__bF_buf10), .S(1'b1) );
DFFSR DFFSR_36 ( .CLK(clk2_clkout_bF_buf5), .D(asr1_rom_2__3_), .Q(asr1_rom_3__3_), .R(_0__bF_buf1), .S(1'b1) );
DFFSR DFFSR_37 ( .CLK(clk2_clkout_bF_buf19), .D(asr1_rom_2__4_), .Q(asr1_rom_3__4_), .R(_0__bF_buf9), .S(1'b1) );
DFFSR DFFSR_38 ( .CLK(clk2_clkout_bF_buf33), .D(asr1_rom_2__5_), .Q(asr1_rom_3__5_), .R(_0__bF_buf5), .S(1'b1) );
DFFSR DFFSR_39 ( .CLK(clk2_clkout_bF_buf34), .D(asr1_rom_2__6_), .Q(asr1_rom_3__6_), .R(_0__bF_buf7), .S(1'b1) );
DFFSR DFFSR_40 ( .CLK(clk2_clkout_bF_buf29), .D(asr1_rom_2__7_), .Q(asr1_rom_3__7_), .R(_0__bF_buf5), .S(1'b1) );
DFFSR DFFSR_41 ( .CLK(clk2_clkout_bF_buf35), .D(asr1_rom_3__0_), .Q(asr1_rom_4__0_), .R(_0__bF_buf9), .S(1'b1) );
DFFSR DFFSR_42 ( .CLK(clk2_clkout_bF_buf33), .D(asr1_rom_3__1_), .Q(asr1_rom_4__1_), .R(_0__bF_buf4), .S(1'b1) );
DFFSR DFFSR_43 ( .CLK(clk2_clkout_bF_buf26), .D(asr1_rom_3__2_), .Q(asr1_rom_4__2_), .R(_0__bF_buf4), .S(1'b1) );
DFFSR DFFSR_44 ( .CLK(clk2_clkout_bF_buf5), .D(asr1_rom_3__3_), .Q(asr1_rom_4__3_), .R(_0__bF_buf1), .S(1'b1) );
DFFSR DFFSR_45 ( .CLK(clk2_clkout_bF_buf0), .D(asr1_rom_3__4_), .Q(asr1_rom_4__4_), .R(_0__bF_buf10), .S(1'b1) );
DFFSR DFFSR_46 ( .CLK(clk2_clkout_bF_buf10), .D(asr1_rom_3__5_), .Q(asr1_rom_4__5_), .R(_0__bF_buf8), .S(1'b1) );
DFFSR DFFSR_47 ( .CLK(clk2_clkout_bF_buf4), .D(asr1_rom_3__6_), .Q(asr1_rom_4__6_), .R(_0__bF_buf6), .S(1'b1) );
DFFSR DFFSR_48 ( .CLK(clk2_clkout_bF_buf29), .D(asr1_rom_3__7_), .Q(asr1_rom_4__7_), .R(_0__bF_buf1), .S(1'b1) );
DFFSR DFFSR_49 ( .CLK(clk2_clkout_bF_buf16), .D(asr1_rom_5__0_), .Q(asr1_rom_6__0_), .R(_0__bF_buf2), .S(1'b1) );
DFFSR DFFSR_50 ( .CLK(clk2_clkout_bF_buf5), .D(asr1_rom_5__1_), .Q(asr1_rom_6__1_), .R(_0__bF_buf1), .S(1'b1) );
DFFSR DFFSR_51 ( .CLK(clk2_clkout_bF_buf34), .D(asr1_rom_5__2_), .Q(asr1_rom_6__2_), .R(_0__bF_buf8), .S(1'b1) );
DFFSR DFFSR_52 ( .CLK(clk2_clkout_bF_buf38), .D(asr1_rom_5__3_), .Q(asr1_rom_6__3_), .R(_0__bF_buf1), .S(1'b1) );
DFFSR DFFSR_53 ( .CLK(clk2_clkout_bF_buf16), .D(asr1_rom_5__4_), .Q(asr1_rom_6__4_), .R(_0__bF_buf2), .S(1'b1) );
DFFSR DFFSR_54 ( .CLK(clk2_clkout_bF_buf10), .D(asr1_rom_5__5_), .Q(asr1_rom_6__5_), .R(_0__bF_buf8), .S(1'b1) );
DFFSR DFFSR_55 ( .CLK(clk2_clkout_bF_buf5), .D(asr1_rom_5__6_), .Q(asr1_rom_6__6_), .R(_0__bF_buf6), .S(1'b1) );
DFFSR DFFSR_56 ( .CLK(clk2_clkout_bF_buf33), .D(asr1_rom_5__7_), .Q(asr1_rom_6__7_), .R(_0__bF_buf4), .S(1'b1) );
DFFSR DFFSR_57 ( .CLK(clk2_clkout_bF_buf26), .D(asr1_rom_4__0_), .Q(asr1_rom_5__0_), .R(_0__bF_buf9), .S(1'b1) );
DFFSR DFFSR_58 ( .CLK(clk2_clkout_bF_buf29), .D(asr1_rom_4__1_), .Q(asr1_rom_5__1_), .R(_0__bF_buf5), .S(1'b1) );
DFFSR DFFSR_59 ( .CLK(clk2_clkout_bF_buf24), .D(asr1_rom_4__2_), .Q(asr1_rom_5__2_), .R(_0__bF_buf3), .S(1'b1) );
DFFSR DFFSR_60 ( .CLK(clk2_clkout_bF_buf38), .D(asr1_rom_4__3_), .Q(asr1_rom_5__3_), .R(_0__bF_buf1), .S(1'b1) );
DFFSR DFFSR_61 ( .CLK(clk2_clkout_bF_buf26), .D(asr1_rom_4__4_), .Q(asr1_rom_5__4_), .R(_0__bF_buf10), .S(1'b1) );
DFFSR DFFSR_62 ( .CLK(clk2_clkout_bF_buf11), .D(asr1_rom_4__5_), .Q(asr1_rom_5__5_), .R(_0__bF_buf8), .S(1'b1) );
DFFSR DFFSR_63 ( .CLK(clk2_clkout_bF_buf4), .D(asr1_rom_4__6_), .Q(asr1_rom_5__6_), .R(_0__bF_buf6), .S(1'b1) );
DFFSR DFFSR_64 ( .CLK(clk2_clkout_bF_buf5), .D(asr1_rom_4__7_), .Q(asr1_rom_5__7_), .R(_0__bF_buf1), .S(1'b1) );
DFFSR DFFSR_65 ( .CLK(clk2_clkout_bF_buf37), .D(asr1_rom_7__0_), .Q(asr1_rom_8__0_), .R(_0__bF_buf4), .S(1'b1) );
DFFSR DFFSR_66 ( .CLK(clk2_clkout_bF_buf7), .D(asr1_rom_7__1_), .Q(asr1_rom_8__1_), .R(_0__bF_buf6), .S(1'b1) );
DFFSR DFFSR_67 ( .CLK(clk2_clkout_bF_buf23), .D(asr1_rom_7__2_), .Q(asr1_rom_8__2_), .R(_0__bF_buf8), .S(1'b1) );
DFFSR DFFSR_68 ( .CLK(clk2_clkout_bF_buf33), .D(asr1_rom_7__3_), .Q(asr1_rom_8__3_), .R(_0__bF_buf4), .S(1'b1) );
DFFSR DFFSR_69 ( .CLK(clk2_clkout_bF_buf26), .D(asr1_rom_7__4_), .Q(asr1_rom_8__4_), .R(_0__bF_buf4), .S(1'b1) );
DFFSR DFFSR_70 ( .CLK(clk2_clkout_bF_buf37), .D(asr1_rom_7__5_), .Q(asr1_rom_8__5_), .R(_0__bF_buf4), .S(1'b1) );
DFFSR DFFSR_71 ( .CLK(clk2_clkout_bF_buf9), .D(asr1_rom_7__6_), .Q(asr1_rom_8__6_), .R(_0__bF_buf7), .S(1'b1) );
DFFSR DFFSR_72 ( .CLK(clk2_clkout_bF_buf37), .D(asr1_rom_7__7_), .Q(asr1_rom_8__7_), .R(_0__bF_buf10), .S(1'b1) );
DFFSR DFFSR_73 ( .CLK(clk2_clkout_bF_buf24), .D(asr1_rom_8__0_), .Q(asr1_rom_9__0_), .R(_0__bF_buf3), .S(1'b1) );
DFFSR DFFSR_74 ( .CLK(clk2_clkout_bF_buf7), .D(asr1_rom_8__1_), .Q(asr1_rom_9__1_), .R(_0__bF_buf10), .S(1'b1) );
DFFSR DFFSR_75 ( .CLK(clk2_clkout_bF_buf10), .D(asr1_rom_8__2_), .Q(asr1_rom_9__2_), .R(_0__bF_buf8), .S(1'b1) );
DFFSR DFFSR_76 ( .CLK(clk2_clkout_bF_buf1), .D(asr1_rom_8__3_), .Q(asr1_rom_9__3_), .R(_0__bF_buf5), .S(1'b1) );
DFFSR DFFSR_77 ( .CLK(clk2_clkout_bF_buf35), .D(asr1_rom_8__4_), .Q(asr1_rom_9__4_), .R(_0__bF_buf9), .S(1'b1) );
DFFSR DFFSR_78 ( .CLK(clk2_clkout_bF_buf0), .D(asr1_rom_8__5_), .Q(asr1_rom_9__5_), .R(_0__bF_buf6), .S(1'b1) );
DFFSR DFFSR_79 ( .CLK(clk2_clkout_bF_buf9), .D(asr1_rom_8__6_), .Q(asr1_rom_9__6_), .R(_0__bF_buf7), .S(1'b1) );
DFFSR DFFSR_80 ( .CLK(clk2_clkout_bF_buf0), .D(asr1_rom_8__7_), .Q(asr1_rom_9__7_), .R(_0__bF_buf10), .S(1'b1) );
DFFSR DFFSR_81 ( .CLK(clk2_clkout_bF_buf34), .D(asr1_rom_9__0_), .Q(asr1_rom_10__0_), .R(_0__bF_buf8), .S(1'b1) );
DFFSR DFFSR_82 ( .CLK(clk2_clkout_bF_buf7), .D(asr1_rom_9__1_), .Q(asr1_rom_10__1_), .R(_0__bF_buf10), .S(1'b1) );
DFFSR DFFSR_83 ( .CLK(clk2_clkout_bF_buf6), .D(asr1_rom_9__2_), .Q(asr1_rom_10__2_), .R(_0__bF_buf3), .S(1'b1) );
DFFSR DFFSR_84 ( .CLK(clk2_clkout_bF_buf1), .D(asr1_rom_9__3_), .Q(asr1_rom_10__3_), .R(_0__bF_buf7), .S(1'b1) );
DFFSR DFFSR_85 ( .CLK(clk2_clkout_bF_buf19), .D(asr1_rom_9__4_), .Q(asr1_rom_10__4_), .R(_0__bF_buf9), .S(1'b1) );
DFFSR DFFSR_86 ( .CLK(clk2_clkout_bF_buf0), .D(asr1_rom_9__5_), .Q(asr1_rom_10__5_), .R(_0__bF_buf6), .S(1'b1) );
DFFSR DFFSR_87 ( .CLK(clk2_clkout_bF_buf4), .D(asr1_rom_9__6_), .Q(asr1_rom_10__6_), .R(_0__bF_buf6), .S(1'b1) );
DFFSR DFFSR_88 ( .CLK(clk2_clkout_bF_buf19), .D(asr1_rom_9__7_), .Q(asr1_rom_10__7_), .R(_0__bF_buf0), .S(1'b1) );
DFFSR DFFSR_89 ( .CLK(clk2_clkout_bF_buf24), .D(asr1_rom_10__0_), .Q(asr1_rom_11__0_), .R(_0__bF_buf3), .S(1'b1) );
DFFSR DFFSR_90 ( .CLK(clk2_clkout_bF_buf7), .D(asr1_rom_10__1_), .Q(asr1_rom_11__1_), .R(_0__bF_buf10), .S(1'b1) );
DFFSR DFFSR_91 ( .CLK(clk2_clkout_bF_buf6), .D(asr1_rom_10__2_), .Q(asr1_rom_11__2_), .R(_0__bF_buf3), .S(1'b1) );
DFFSR DFFSR_92 ( .CLK(clk2_clkout_bF_buf1), .D(asr1_rom_10__3_), .Q(asr1_rom_11__3_), .R(_0__bF_buf7), .S(1'b1) );
DFFSR DFFSR_93 ( .CLK(clk2_clkout_bF_buf18), .D(asr1_rom_10__4_), .Q(asr1_rom_11__4_), .R(_0__bF_buf0), .S(1'b1) );
DFFSR DFFSR_94 ( .CLK(clk2_clkout_bF_buf4), .D(asr1_rom_10__5_), .Q(asr1_rom_11__5_), .R(_0__bF_buf6), .S(1'b1) );
DFFSR DFFSR_95 ( .CLK(clk2_clkout_bF_buf4), .D(asr1_rom_10__6_), .Q(asr1_rom_11__6_), .R(_0__bF_buf6), .S(1'b1) );
DFFSR DFFSR_96 ( .CLK(clk2_clkout_bF_buf19), .D(asr1_rom_10__7_), .Q(asr1_rom_11__7_), .R(_0__bF_buf0), .S(1'b1) );
DFFSR DFFSR_97 ( .CLK(clk2_clkout_bF_buf6), .D(asr1_rom_11__0_), .Q(asr1_rom_12__0_), .R(_0__bF_buf3), .S(1'b1) );
DFFSR DFFSR_98 ( .CLK(clk2_clkout_bF_buf7), .D(asr1_rom_11__1_), .Q(asr1_rom_12__1_), .R(_0__bF_buf0), .S(1'b1) );
DFFSR DFFSR_99 ( .CLK(clk2_clkout_bF_buf6), .D(asr1_rom_11__2_), .Q(asr1_rom_12__2_), .R(_0__bF_buf3), .S(1'b1) );
DFFSR DFFSR_100 ( .CLK(clk2_clkout_bF_buf9), .D(asr1_rom_11__3_), .Q(asr1_rom_12__3_), .R(_0__bF_buf7), .S(1'b1) );
DFFSR DFFSR_101 ( .CLK(clk2_clkout_bF_buf18), .D(asr1_rom_11__4_), .Q(asr1_rom_12__4_), .R(_0__bF_buf0), .S(1'b1) );
DFFSR DFFSR_102 ( .CLK(clk2_clkout_bF_buf0), .D(asr1_rom_11__5_), .Q(asr1_rom_12__5_), .R(_0__bF_buf6), .S(1'b1) );
DFFSR DFFSR_103 ( .CLK(clk2_clkout_bF_buf37), .D(asr1_rom_11__6_), .Q(asr1_rom_12__6_), .R(_0__bF_buf4), .S(1'b1) );
DFFSR DFFSR_104 ( .CLK(clk2_clkout_bF_buf35), .D(asr1_rom_11__7_), .Q(asr1_rom_12__7_), .R(_0__bF_buf10), .S(1'b1) );
DFFSR DFFSR_105 ( .CLK(clk2_clkout_bF_buf16), .D(asr1_rom_12__0_), .Q(asr1_rom_13__0_), .R(_0__bF_buf2), .S(1'b1) );
DFFSR DFFSR_106 ( .CLK(clk2_clkout_bF_buf15), .D(asr1_rom_12__1_), .Q(asr1_rom_13__1_), .R(_0__bF_buf2), .S(1'b1) );
DFFSR DFFSR_107 ( .CLK(clk2_clkout_bF_buf16), .D(asr1_rom_12__2_), .Q(asr1_rom_13__2_), .R(_0__bF_buf3), .S(1'b1) );
DFFSR DFFSR_108 ( .CLK(clk2_clkout_bF_buf9), .D(asr1_rom_12__3_), .Q(asr1_rom_13__3_), .R(_0__bF_buf7), .S(1'b1) );
DFFSR DFFSR_109 ( .CLK(clk2_clkout_bF_buf18), .D(asr1_rom_12__4_), .Q(asr1_rom_13__4_), .R(_0__bF_buf0), .S(1'b1) );
DFFSR DFFSR_110 ( .CLK(clk2_clkout_bF_buf0), .D(asr1_rom_12__5_), .Q(asr1_rom_13__5_), .R(_0__bF_buf10), .S(1'b1) );
DFFSR DFFSR_111 ( .CLK(clk2_clkout_bF_buf37), .D(asr1_rom_12__6_), .Q(asr1_rom_13__6_), .R(_0__bF_buf10), .S(1'b1) );
DFFSR DFFSR_112 ( .CLK(clk2_clkout_bF_buf26), .D(asr1_rom_12__7_), .Q(asr1_rom_13__7_), .R(_0__bF_buf9), .S(1'b1) );
DFFSR DFFSR_113 ( .CLK(clk2_clkout_bF_buf2), .D(asr1_rom_13__0_), .Q(asr1_rom_14__0_), .R(_0__bF_buf2), .S(1'b1) );
DFFSR DFFSR_114 ( .CLK(clk2_clkout_bF_buf15), .D(asr1_rom_13__1_), .Q(asr1_rom_14__1_), .R(_0__bF_buf2), .S(1'b1) );
DFFSR DFFSR_115 ( .CLK(clk2_clkout_bF_buf15), .D(asr1_rom_13__2_), .Q(asr1_rom_14__2_), .R(_0__bF_buf2), .S(1'b1) );
DFFSR DFFSR_116 ( .CLK(clk2_clkout_bF_buf34), .D(asr1_rom_13__3_), .Q(asr1_rom_14__3_), .R(_0__bF_buf7), .S(1'b1) );
DFFSR DFFSR_117 ( .CLK(clk2_clkout_bF_buf18), .D(asr1_rom_13__4_), .Q(asr1_rom_14__4_), .R(_0__bF_buf0), .S(1'b1) );
DFFSR DFFSR_118 ( .CLK(clk2_clkout_bF_buf26), .D(asr1_rom_13__5_), .Q(asr1_rom_14__5_), .R(_0__bF_buf10), .S(1'b1) );
DFFSR DFFSR_119 ( .CLK(clk2_clkout_bF_buf37), .D(asr1_rom_13__6_), .Q(asr1_rom_14__6_), .R(_0__bF_buf4), .S(1'b1) );
DFFSR DFFSR_120 ( .CLK(clk2_clkout_bF_buf24), .D(asr1_rom_13__7_), .Q(asr1_rom_14__7_), .R(_0__bF_buf3), .S(1'b1) );
DFFSR DFFSR_121 ( .CLK(clk2_clkout_bF_buf2), .D(asr1_rom_14__0_), .Q(asr1_en_0_), .R(_0__bF_buf2), .S(1'b1) );
DFFSR DFFSR_122 ( .CLK(clk2_clkout_bF_buf2), .D(asr1_rom_14__1_), .Q(asr1_en_1_), .R(_0__bF_buf2), .S(1'b1) );
DFFSR DFFSR_123 ( .CLK(clk2_clkout_bF_buf15), .D(asr1_rom_14__2_), .Q(asr1_en_2_), .R(_0__bF_buf2), .S(1'b1) );
DFFSR DFFSR_124 ( .CLK(clk2_clkout_bF_buf34), .D(asr1_rom_14__3_), .Q(asr1_en_3_), .R(_0__bF_buf8), .S(1'b1) );
DFFSR DFFSR_125 ( .CLK(clk2_clkout_bF_buf18), .D(asr1_rom_14__4_), .Q(asr1_en_4_), .R(_0__bF_buf0), .S(1'b1) );
DFFSR DFFSR_126 ( .CLK(clk2_clkout_bF_buf2), .D(asr1_rom_14__5_), .Q(asr1_en_5_), .R(_0__bF_buf2), .S(1'b1) );
DFFSR DFFSR_127 ( .CLK(clk2_clkout_bF_buf37), .D(asr1_rom_14__6_), .Q(asr1_en_6_), .R(_0__bF_buf7), .S(1'b1) );
DFFSR DFFSR_128 ( .CLK(clk2_clkout_bF_buf6), .D(asr1_rom_14__7_), .Q(asr1_en_7_), .R(_0__bF_buf3), .S(1'b1) );
INVX1 INVX1_60 ( .A(asr2_rom_6__0_), .Y(_226_) );
INVX1 INVX1_61 ( .A(asr2_rom_5__0_), .Y(_227_) );
INVX1 INVX1_62 ( .A(counterdown_counter_3_), .Y(_228_) );
AND2X2 AND2X2_14 ( .A(_228_), .B(counterdown_counter_2_), .Y(_229_) );
INVX1 INVX1_63 ( .A(counterdown_counter_1_), .Y(_230_) );
AND2X2 AND2X2_15 ( .A(_230_), .B(counterdown_counter_0_), .Y(_231_) );
NAND2X1 NAND2X1_27 ( .A(_229__bF_buf1), .B(_231_), .Y(_232_) );
NOR2X1 NOR2X1_30 ( .A(counterdown_counter_0_), .B(_230_), .Y(_233_) );
NAND2X1 NAND2X1_28 ( .A(_233_), .B(_229__bF_buf1), .Y(_234_) );
OAI22X1 OAI22X1_25 ( .A(_226_), .B(_234_), .C(_227_), .D(_232_), .Y(_235_) );
INVX1 INVX1_64 ( .A(asr2_rom_10__0_), .Y(_236_) );
INVX1 INVX1_65 ( .A(asr2_rom_9__0_), .Y(_237_) );
NOR2X1 NOR2X1_31 ( .A(counterdown_counter_2_), .B(_228_), .Y(_238_) );
NAND2X1 NAND2X1_29 ( .A(_238_), .B(_231_), .Y(_239_) );
NAND2X1 NAND2X1_30 ( .A(_233_), .B(_238_), .Y(_240_) );
OAI22X1 OAI22X1_26 ( .A(_236_), .B(_240_), .C(_237_), .D(_239_), .Y(_241_) );
NOR2X1 NOR2X1_32 ( .A(_241_), .B(_235_), .Y(_242_) );
INVX1 INVX1_66 ( .A(asr2_rom_2__0_), .Y(_243_) );
INVX1 INVX1_67 ( .A(asr2_rom_1__0_), .Y(_244_) );
NOR2X1 NOR2X1_33 ( .A(counterdown_counter_3_), .B(counterdown_counter_2_), .Y(_245_) );
NAND2X1 NAND2X1_31 ( .A(_245_), .B(_231_), .Y(_246_) );
NAND2X1 NAND2X1_32 ( .A(_245_), .B(_233_), .Y(_247_) );
OAI22X1 OAI22X1_27 ( .A(_243_), .B(_247_), .C(_244_), .D(_246_), .Y(_248_) );
INVX1 INVX1_68 ( .A(asr2_rom_14__0_), .Y(_249_) );
NAND2X1 NAND2X1_33 ( .A(counterdown_counter_0_), .B(_230_), .Y(_250_) );
NAND2X1 NAND2X1_34 ( .A(counterdown_counter_3_), .B(counterdown_counter_2_), .Y(_251_) );
NOR2X1 NOR2X1_34 ( .A(_251_), .B(_250_), .Y(_252_) );
NAND2X1 NAND2X1_35 ( .A(asr2_rom_13__0_), .B(_252_), .Y(_253_) );
AND2X2 AND2X2_16 ( .A(counterdown_counter_3_), .B(counterdown_counter_2_), .Y(_254_) );
NAND2X1 NAND2X1_36 ( .A(_254_), .B(_233_), .Y(_255_) );
OAI21X1 OAI21X1_9 ( .A(_249_), .B(_255_), .C(_253_), .Y(_256_) );
NOR2X1 NOR2X1_35 ( .A(_248_), .B(_256_), .Y(_257_) );
AND2X2 AND2X2_17 ( .A(counterdown_counter_1_), .B(counterdown_counter_0_), .Y(_258_) );
AND2X2 AND2X2_18 ( .A(_258__bF_buf2), .B(_245_), .Y(_259_) );
NAND2X1 NAND2X1_37 ( .A(asr2_rom_3__0_), .B(_259_), .Y(_260_) );
NOR2X1 NOR2X1_36 ( .A(counterdown_counter_1_), .B(counterdown_counter_0_), .Y(_261_) );
NAND3X1 NAND3X1_65 ( .A(asr2_rom_4__0_), .B(_261__bF_buf3), .C(_229__bF_buf3), .Y(_262_) );
NAND3X1 NAND3X1_66 ( .A(asr2_rom_0__0_), .B(_245_), .C(_261__bF_buf3), .Y(_263_) );
NAND3X1 NAND3X1_67 ( .A(asr2_en_0_), .B(_254_), .C(_258__bF_buf0), .Y(_264_) );
AND2X2 AND2X2_19 ( .A(_264_), .B(_263_), .Y(_265_) );
NAND3X1 NAND3X1_68 ( .A(_260_), .B(_262_), .C(_265_), .Y(_266_) );
NAND3X1 NAND3X1_69 ( .A(asr2_rom_7__0_), .B(_258__bF_buf3), .C(_229__bF_buf2), .Y(_267_) );
NAND3X1 NAND3X1_70 ( .A(asr2_rom_8__0_), .B(_261__bF_buf2), .C(_238_), .Y(_268_) );
NAND2X1 NAND2X1_38 ( .A(counterdown_counter_1_), .B(counterdown_counter_0_), .Y(_269_) );
NOR3X1 NOR3X1_3 ( .A(counterdown_counter_2_), .B(_228_), .C(_269_), .Y(_270_) );
NOR3X1 NOR3X1_4 ( .A(counterdown_counter_1_), .B(counterdown_counter_0_), .C(_251_), .Y(_271_) );
AOI22X1 AOI22X1_9 ( .A(_271_), .B(asr2_rom_12__0_), .C(asr2_rom_11__0_), .D(_270_), .Y(_272_) );
NAND3X1 NAND3X1_71 ( .A(_267_), .B(_268_), .C(_272_), .Y(_273_) );
NOR2X1 NOR2X1_37 ( .A(_266_), .B(_273_), .Y(_274_) );
NAND3X1 NAND3X1_72 ( .A(_242_), .B(_257_), .C(_274_), .Y(asr2_dataout_0_) );
INVX1 INVX1_69 ( .A(asr2_rom_6__1_), .Y(_275_) );
INVX1 INVX1_70 ( .A(asr2_rom_5__1_), .Y(_276_) );
OAI22X1 OAI22X1_28 ( .A(_275_), .B(_234_), .C(_276_), .D(_232_), .Y(_277_) );
INVX1 INVX1_71 ( .A(asr2_rom_10__1_), .Y(_278_) );
INVX1 INVX1_72 ( .A(asr2_rom_9__1_), .Y(_279_) );
OAI22X1 OAI22X1_29 ( .A(_278_), .B(_240_), .C(_279_), .D(_239_), .Y(_280_) );
NOR2X1 NOR2X1_38 ( .A(_280_), .B(_277_), .Y(_281_) );
INVX1 INVX1_73 ( .A(asr2_rom_2__1_), .Y(_282_) );
INVX1 INVX1_74 ( .A(asr2_rom_1__1_), .Y(_283_) );
OAI22X1 OAI22X1_30 ( .A(_282_), .B(_247_), .C(_283_), .D(_246_), .Y(_284_) );
INVX1 INVX1_75 ( .A(asr2_rom_14__1_), .Y(_285_) );
NAND2X1 NAND2X1_39 ( .A(asr2_rom_13__1_), .B(_252_), .Y(_286_) );
OAI21X1 OAI21X1_10 ( .A(_285_), .B(_255_), .C(_286_), .Y(_287_) );
NOR2X1 NOR2X1_39 ( .A(_284_), .B(_287_), .Y(_288_) );
NAND2X1 NAND2X1_40 ( .A(asr2_rom_3__1_), .B(_259_), .Y(_289_) );
NAND3X1 NAND3X1_73 ( .A(asr2_rom_4__1_), .B(_261__bF_buf0), .C(_229__bF_buf0), .Y(_290_) );
NAND3X1 NAND3X1_74 ( .A(asr2_rom_0__1_), .B(_245_), .C(_261__bF_buf0), .Y(_291_) );
NAND3X1 NAND3X1_75 ( .A(asr2_en_1_), .B(_254_), .C(_258__bF_buf1), .Y(_292_) );
AND2X2 AND2X2_20 ( .A(_292_), .B(_291_), .Y(_293_) );
NAND3X1 NAND3X1_76 ( .A(_289_), .B(_290_), .C(_293_), .Y(_294_) );
NAND3X1 NAND3X1_77 ( .A(asr2_rom_7__1_), .B(_258__bF_buf3), .C(_229__bF_buf2), .Y(_295_) );
NAND3X1 NAND3X1_78 ( .A(asr2_rom_8__1_), .B(_261__bF_buf0), .C(_238_), .Y(_296_) );
AOI22X1 AOI22X1_10 ( .A(_271_), .B(asr2_rom_12__1_), .C(asr2_rom_11__1_), .D(_270_), .Y(_297_) );
NAND3X1 NAND3X1_79 ( .A(_295_), .B(_296_), .C(_297_), .Y(_298_) );
NOR2X1 NOR2X1_40 ( .A(_294_), .B(_298_), .Y(_299_) );
NAND3X1 NAND3X1_80 ( .A(_281_), .B(_288_), .C(_299_), .Y(asr2_dataout_1_) );
INVX1 INVX1_76 ( .A(asr2_rom_6__2_), .Y(_300_) );
INVX1 INVX1_77 ( .A(asr2_rom_5__2_), .Y(_301_) );
OAI22X1 OAI22X1_31 ( .A(_300_), .B(_234_), .C(_301_), .D(_232_), .Y(_302_) );
INVX1 INVX1_78 ( .A(asr2_rom_10__2_), .Y(_303_) );
INVX1 INVX1_79 ( .A(asr2_rom_9__2_), .Y(_304_) );
OAI22X1 OAI22X1_32 ( .A(_303_), .B(_240_), .C(_304_), .D(_239_), .Y(_305_) );
NOR2X1 NOR2X1_41 ( .A(_305_), .B(_302_), .Y(_306_) );
INVX1 INVX1_80 ( .A(asr2_rom_2__2_), .Y(_307_) );
INVX1 INVX1_81 ( .A(asr2_rom_1__2_), .Y(_308_) );
OAI22X1 OAI22X1_33 ( .A(_307_), .B(_247_), .C(_308_), .D(_246_), .Y(_309_) );
INVX1 INVX1_82 ( .A(asr2_rom_14__2_), .Y(_310_) );
NAND2X1 NAND2X1_41 ( .A(asr2_rom_13__2_), .B(_252_), .Y(_311_) );
OAI21X1 OAI21X1_11 ( .A(_310_), .B(_255_), .C(_311_), .Y(_312_) );
NOR2X1 NOR2X1_42 ( .A(_309_), .B(_312_), .Y(_313_) );
NAND2X1 NAND2X1_42 ( .A(asr2_rom_3__2_), .B(_259_), .Y(_314_) );
NAND3X1 NAND3X1_81 ( .A(asr2_rom_4__2_), .B(_261__bF_buf1), .C(_229__bF_buf1), .Y(_315_) );
NAND3X1 NAND3X1_82 ( .A(asr2_rom_0__2_), .B(_245_), .C(_261__bF_buf2), .Y(_316_) );
NAND3X1 NAND3X1_83 ( .A(asr2_en_2_), .B(_254_), .C(_258__bF_buf3), .Y(_317_) );
AND2X2 AND2X2_21 ( .A(_317_), .B(_316_), .Y(_318_) );
NAND3X1 NAND3X1_84 ( .A(_314_), .B(_315_), .C(_318_), .Y(_319_) );
NAND3X1 NAND3X1_85 ( .A(asr2_rom_7__2_), .B(_258__bF_buf0), .C(_229__bF_buf3), .Y(_320_) );
NAND3X1 NAND3X1_86 ( .A(asr2_rom_8__2_), .B(_261__bF_buf3), .C(_238_), .Y(_321_) );
AOI22X1 AOI22X1_11 ( .A(_271_), .B(asr2_rom_12__2_), .C(asr2_rom_11__2_), .D(_270_), .Y(_322_) );
NAND3X1 NAND3X1_87 ( .A(_320_), .B(_321_), .C(_322_), .Y(_323_) );
NOR2X1 NOR2X1_43 ( .A(_319_), .B(_323_), .Y(_324_) );
NAND3X1 NAND3X1_88 ( .A(_306_), .B(_313_), .C(_324_), .Y(asr2_dataout_2_) );
INVX1 INVX1_83 ( .A(asr2_rom_6__3_), .Y(_325_) );
INVX1 INVX1_84 ( .A(asr2_rom_5__3_), .Y(_326_) );
OAI22X1 OAI22X1_34 ( .A(_325_), .B(_234_), .C(_326_), .D(_232_), .Y(_327_) );
INVX1 INVX1_85 ( .A(asr2_rom_10__3_), .Y(_328_) );
INVX1 INVX1_86 ( .A(asr2_rom_9__3_), .Y(_329_) );
OAI22X1 OAI22X1_35 ( .A(_328_), .B(_240_), .C(_329_), .D(_239_), .Y(_330_) );
NOR2X1 NOR2X1_44 ( .A(_330_), .B(_327_), .Y(_331_) );
INVX1 INVX1_87 ( .A(asr2_rom_2__3_), .Y(_332_) );
INVX1 INVX1_88 ( .A(asr2_rom_1__3_), .Y(_333_) );
OAI22X1 OAI22X1_36 ( .A(_332_), .B(_247_), .C(_333_), .D(_246_), .Y(_334_) );
INVX1 INVX1_89 ( .A(asr2_rom_14__3_), .Y(_335_) );
NAND2X1 NAND2X1_43 ( .A(asr2_rom_13__3_), .B(_252_), .Y(_336_) );
OAI21X1 OAI21X1_12 ( .A(_335_), .B(_255_), .C(_336_), .Y(_337_) );
NOR2X1 NOR2X1_45 ( .A(_334_), .B(_337_), .Y(_338_) );
NAND2X1 NAND2X1_44 ( .A(asr2_rom_3__3_), .B(_259_), .Y(_339_) );
NAND3X1 NAND3X1_89 ( .A(asr2_rom_4__3_), .B(_261__bF_buf3), .C(_229__bF_buf3), .Y(_340_) );
NAND3X1 NAND3X1_90 ( .A(asr2_rom_0__3_), .B(_245_), .C(_261__bF_buf1), .Y(_341_) );
NAND3X1 NAND3X1_91 ( .A(asr2_en_3_), .B(_254_), .C(_258__bF_buf2), .Y(_342_) );
AND2X2 AND2X2_22 ( .A(_342_), .B(_341_), .Y(_343_) );
NAND3X1 NAND3X1_92 ( .A(_339_), .B(_340_), .C(_343_), .Y(_344_) );
NAND3X1 NAND3X1_93 ( .A(asr2_rom_7__3_), .B(_258__bF_buf0), .C(_229__bF_buf3), .Y(_345_) );
NAND3X1 NAND3X1_94 ( .A(asr2_rom_8__3_), .B(_261__bF_buf3), .C(_238_), .Y(_346_) );
AOI22X1 AOI22X1_12 ( .A(_271_), .B(asr2_rom_12__3_), .C(asr2_rom_11__3_), .D(_270_), .Y(_347_) );
NAND3X1 NAND3X1_95 ( .A(_345_), .B(_346_), .C(_347_), .Y(_348_) );
NOR2X1 NOR2X1_46 ( .A(_344_), .B(_348_), .Y(_349_) );
NAND3X1 NAND3X1_96 ( .A(_331_), .B(_338_), .C(_349_), .Y(asr2_dataout_3_) );
INVX1 INVX1_90 ( .A(asr2_rom_6__4_), .Y(_350_) );
INVX1 INVX1_91 ( .A(asr2_rom_5__4_), .Y(_351_) );
OAI22X1 OAI22X1_37 ( .A(_350_), .B(_234_), .C(_351_), .D(_232_), .Y(_352_) );
INVX1 INVX1_92 ( .A(asr2_rom_10__4_), .Y(_353_) );
INVX1 INVX1_93 ( .A(asr2_rom_9__4_), .Y(_354_) );
OAI22X1 OAI22X1_38 ( .A(_353_), .B(_240_), .C(_354_), .D(_239_), .Y(_355_) );
NOR2X1 NOR2X1_47 ( .A(_355_), .B(_352_), .Y(_356_) );
INVX1 INVX1_94 ( .A(asr2_rom_2__4_), .Y(_357_) );
INVX1 INVX1_95 ( .A(asr2_rom_1__4_), .Y(_358_) );
OAI22X1 OAI22X1_39 ( .A(_357_), .B(_247_), .C(_358_), .D(_246_), .Y(_359_) );
INVX1 INVX1_96 ( .A(asr2_rom_14__4_), .Y(_360_) );
NAND2X1 NAND2X1_45 ( .A(asr2_rom_13__4_), .B(_252_), .Y(_361_) );
OAI21X1 OAI21X1_13 ( .A(_360_), .B(_255_), .C(_361_), .Y(_362_) );
NOR2X1 NOR2X1_48 ( .A(_359_), .B(_362_), .Y(_363_) );
NAND2X1 NAND2X1_46 ( .A(asr2_rom_3__4_), .B(_259_), .Y(_364_) );
NAND3X1 NAND3X1_97 ( .A(asr2_rom_4__4_), .B(_261__bF_buf0), .C(_229__bF_buf0), .Y(_365_) );
NAND3X1 NAND3X1_98 ( .A(asr2_rom_0__4_), .B(_245_), .C(_261__bF_buf1), .Y(_366_) );
NAND3X1 NAND3X1_99 ( .A(asr2_en_4_), .B(_254_), .C(_258__bF_buf2), .Y(_367_) );
AND2X2 AND2X2_23 ( .A(_367_), .B(_366_), .Y(_368_) );
NAND3X1 NAND3X1_100 ( .A(_364_), .B(_365_), .C(_368_), .Y(_369_) );
NAND3X1 NAND3X1_101 ( .A(asr2_rom_7__4_), .B(_258__bF_buf1), .C(_229__bF_buf0), .Y(_370_) );
NAND3X1 NAND3X1_102 ( .A(asr2_rom_8__4_), .B(_261__bF_buf1), .C(_238_), .Y(_371_) );
AOI22X1 AOI22X1_13 ( .A(_271_), .B(asr2_rom_12__4_), .C(asr2_rom_11__4_), .D(_270_), .Y(_372_) );
NAND3X1 NAND3X1_103 ( .A(_370_), .B(_371_), .C(_372_), .Y(_373_) );
NOR2X1 NOR2X1_49 ( .A(_369_), .B(_373_), .Y(_374_) );
NAND3X1 NAND3X1_104 ( .A(_356_), .B(_363_), .C(_374_), .Y(asr2_dataout_4_) );
INVX1 INVX1_97 ( .A(asr2_rom_6__5_), .Y(_375_) );
INVX1 INVX1_98 ( .A(asr2_rom_5__5_), .Y(_376_) );
OAI22X1 OAI22X1_40 ( .A(_375_), .B(_234_), .C(_376_), .D(_232_), .Y(_377_) );
INVX1 INVX1_99 ( .A(asr2_rom_10__5_), .Y(_378_) );
INVX1 INVX1_100 ( .A(asr2_rom_9__5_), .Y(_379_) );
OAI22X1 OAI22X1_41 ( .A(_378_), .B(_240_), .C(_379_), .D(_239_), .Y(_380_) );
NOR2X1 NOR2X1_50 ( .A(_380_), .B(_377_), .Y(_381_) );
INVX1 INVX1_101 ( .A(asr2_rom_2__5_), .Y(_382_) );
INVX1 INVX1_102 ( .A(asr2_rom_1__5_), .Y(_383_) );
OAI22X1 OAI22X1_42 ( .A(_382_), .B(_247_), .C(_383_), .D(_246_), .Y(_384_) );
INVX1 INVX1_103 ( .A(asr2_rom_14__5_), .Y(_385_) );
NAND2X1 NAND2X1_47 ( .A(asr2_rom_13__5_), .B(_252_), .Y(_386_) );
OAI21X1 OAI21X1_14 ( .A(_385_), .B(_255_), .C(_386_), .Y(_387_) );
NOR2X1 NOR2X1_51 ( .A(_384_), .B(_387_), .Y(_388_) );
NAND2X1 NAND2X1_48 ( .A(asr2_rom_3__5_), .B(_259_), .Y(_389_) );
NAND3X1 NAND3X1_105 ( .A(asr2_rom_4__5_), .B(_261__bF_buf1), .C(_229__bF_buf1), .Y(_390_) );
NAND3X1 NAND3X1_106 ( .A(asr2_rom_0__5_), .B(_245_), .C(_261__bF_buf1), .Y(_391_) );
NAND3X1 NAND3X1_107 ( .A(asr2_en_5_), .B(_254_), .C(_258__bF_buf2), .Y(_392_) );
AND2X2 AND2X2_24 ( .A(_392_), .B(_391_), .Y(_393_) );
NAND3X1 NAND3X1_108 ( .A(_389_), .B(_390_), .C(_393_), .Y(_394_) );
NAND3X1 NAND3X1_109 ( .A(asr2_rom_7__5_), .B(_258__bF_buf0), .C(_229__bF_buf3), .Y(_395_) );
NAND3X1 NAND3X1_110 ( .A(asr2_rom_8__5_), .B(_261__bF_buf3), .C(_238_), .Y(_396_) );
AOI22X1 AOI22X1_14 ( .A(_271_), .B(asr2_rom_12__5_), .C(asr2_rom_11__5_), .D(_270_), .Y(_397_) );
NAND3X1 NAND3X1_111 ( .A(_395_), .B(_396_), .C(_397_), .Y(_398_) );
NOR2X1 NOR2X1_52 ( .A(_394_), .B(_398_), .Y(_399_) );
NAND3X1 NAND3X1_112 ( .A(_381_), .B(_388_), .C(_399_), .Y(asr2_dataout_5_) );
INVX1 INVX1_104 ( .A(asr2_rom_6__6_), .Y(_400_) );
INVX1 INVX1_105 ( .A(asr2_rom_5__6_), .Y(_401_) );
OAI22X1 OAI22X1_43 ( .A(_400_), .B(_234_), .C(_401_), .D(_232_), .Y(_402_) );
INVX1 INVX1_106 ( .A(asr2_rom_10__6_), .Y(_403_) );
INVX1 INVX1_107 ( .A(asr2_rom_9__6_), .Y(_404_) );
OAI22X1 OAI22X1_44 ( .A(_403_), .B(_240_), .C(_404_), .D(_239_), .Y(_405_) );
NOR2X1 NOR2X1_53 ( .A(_405_), .B(_402_), .Y(_406_) );
INVX1 INVX1_108 ( .A(asr2_rom_2__6_), .Y(_407_) );
INVX1 INVX1_109 ( .A(asr2_rom_1__6_), .Y(_408_) );
OAI22X1 OAI22X1_45 ( .A(_407_), .B(_247_), .C(_408_), .D(_246_), .Y(_409_) );
INVX1 INVX1_110 ( .A(asr2_rom_14__6_), .Y(_410_) );
NAND2X1 NAND2X1_49 ( .A(asr2_rom_13__6_), .B(_252_), .Y(_411_) );
OAI21X1 OAI21X1_15 ( .A(_410_), .B(_255_), .C(_411_), .Y(_412_) );
NOR2X1 NOR2X1_54 ( .A(_409_), .B(_412_), .Y(_413_) );
NAND2X1 NAND2X1_50 ( .A(asr2_rom_3__6_), .B(_259_), .Y(_414_) );
NAND3X1 NAND3X1_113 ( .A(asr2_rom_4__6_), .B(_261__bF_buf2), .C(_229__bF_buf2), .Y(_415_) );
NAND3X1 NAND3X1_114 ( .A(asr2_rom_0__6_), .B(_245_), .C(_261__bF_buf2), .Y(_416_) );
NAND3X1 NAND3X1_115 ( .A(asr2_en_6_), .B(_254_), .C(_258__bF_buf1), .Y(_417_) );
AND2X2 AND2X2_25 ( .A(_417_), .B(_416_), .Y(_418_) );
NAND3X1 NAND3X1_116 ( .A(_414_), .B(_415_), .C(_418_), .Y(_419_) );
NAND3X1 NAND3X1_117 ( .A(asr2_rom_7__6_), .B(_258__bF_buf3), .C(_229__bF_buf2), .Y(_420_) );
NAND3X1 NAND3X1_118 ( .A(asr2_rom_8__6_), .B(_261__bF_buf2), .C(_238_), .Y(_421_) );
AOI22X1 AOI22X1_15 ( .A(_271_), .B(asr2_rom_12__6_), .C(asr2_rom_11__6_), .D(_270_), .Y(_422_) );
NAND3X1 NAND3X1_119 ( .A(_420_), .B(_421_), .C(_422_), .Y(_423_) );
NOR2X1 NOR2X1_55 ( .A(_419_), .B(_423_), .Y(_424_) );
NAND3X1 NAND3X1_120 ( .A(_406_), .B(_413_), .C(_424_), .Y(asr2_dataout_6_) );
INVX1 INVX1_111 ( .A(asr2_rom_6__7_), .Y(_425_) );
INVX1 INVX1_112 ( .A(asr2_rom_5__7_), .Y(_426_) );
OAI22X1 OAI22X1_46 ( .A(_425_), .B(_234_), .C(_426_), .D(_232_), .Y(_427_) );
INVX1 INVX1_113 ( .A(asr2_rom_10__7_), .Y(_428_) );
INVX1 INVX1_114 ( .A(asr2_rom_9__7_), .Y(_429_) );
OAI22X1 OAI22X1_47 ( .A(_428_), .B(_240_), .C(_429_), .D(_239_), .Y(_430_) );
NOR2X1 NOR2X1_56 ( .A(_430_), .B(_427_), .Y(_431_) );
INVX1 INVX1_115 ( .A(asr2_rom_2__7_), .Y(_432_) );
INVX1 INVX1_116 ( .A(asr2_rom_1__7_), .Y(_433_) );
OAI22X1 OAI22X1_48 ( .A(_432_), .B(_247_), .C(_433_), .D(_246_), .Y(_434_) );
INVX1 INVX1_117 ( .A(asr2_rom_14__7_), .Y(_435_) );
NAND2X1 NAND2X1_51 ( .A(asr2_rom_13__7_), .B(_252_), .Y(_436_) );
OAI21X1 OAI21X1_16 ( .A(_435_), .B(_255_), .C(_436_), .Y(_437_) );
NOR2X1 NOR2X1_57 ( .A(_434_), .B(_437_), .Y(_438_) );
NAND2X1 NAND2X1_52 ( .A(asr2_rom_3__7_), .B(_259_), .Y(_439_) );
NAND3X1 NAND3X1_121 ( .A(asr2_rom_4__7_), .B(_261__bF_buf0), .C(_229__bF_buf0), .Y(_440_) );
NAND3X1 NAND3X1_122 ( .A(asr2_rom_0__7_), .B(_245_), .C(_261__bF_buf0), .Y(_441_) );
NAND3X1 NAND3X1_123 ( .A(asr2_en_7_), .B(_254_), .C(_258__bF_buf1), .Y(_442_) );
AND2X2 AND2X2_26 ( .A(_442_), .B(_441_), .Y(_443_) );
NAND3X1 NAND3X1_124 ( .A(_439_), .B(_440_), .C(_443_), .Y(_444_) );
NAND3X1 NAND3X1_125 ( .A(asr2_rom_7__7_), .B(_258__bF_buf3), .C(_229__bF_buf2), .Y(_445_) );
NAND3X1 NAND3X1_126 ( .A(asr2_rom_8__7_), .B(_261__bF_buf2), .C(_238_), .Y(_446_) );
AOI22X1 AOI22X1_16 ( .A(_271_), .B(asr2_rom_12__7_), .C(asr2_rom_11__7_), .D(_270_), .Y(_447_) );
NAND3X1 NAND3X1_127 ( .A(_445_), .B(_446_), .C(_447_), .Y(_448_) );
NOR2X1 NOR2X1_58 ( .A(_444_), .B(_448_), .Y(_449_) );
NAND3X1 NAND3X1_128 ( .A(_431_), .B(_438_), .C(_449_), .Y(asr2_dataout_7_) );
INVX1 INVX1_118 ( .A(rst_bF_buf0), .Y(_225_) );
DFFSR DFFSR_129 ( .CLK(clk2_clkout_bF_buf31), .D(asr1_en_0_), .Q(asr2_rom_0__0_), .R(_225__bF_buf3), .S(1'b1) );
DFFSR DFFSR_130 ( .CLK(clk2_clkout_bF_buf39), .D(asr1_en_1_), .Q(asr2_rom_0__1_), .R(_225__bF_buf7), .S(1'b1) );
DFFSR DFFSR_131 ( .CLK(clk2_clkout_bF_buf15), .D(asr1_en_2_), .Q(asr2_rom_0__2_), .R(_225__bF_buf9), .S(1'b1) );
DFFSR DFFSR_132 ( .CLK(clk2_clkout_bF_buf24), .D(asr1_en_3_), .Q(asr2_rom_0__3_), .R(_225__bF_buf9), .S(1'b1) );
DFFSR DFFSR_133 ( .CLK(clk2_clkout_bF_buf12), .D(asr1_en_4_), .Q(asr2_rom_0__4_), .R(_225__bF_buf5), .S(1'b1) );
DFFSR DFFSR_134 ( .CLK(clk2_clkout_bF_buf2), .D(asr1_en_5_), .Q(asr2_rom_0__5_), .R(_225__bF_buf7), .S(1'b1) );
DFFSR DFFSR_135 ( .CLK(clk2_clkout_bF_buf11), .D(asr1_en_6_), .Q(asr2_rom_0__6_), .R(_225__bF_buf2), .S(1'b1) );
DFFSR DFFSR_136 ( .CLK(clk2_clkout_bF_buf15), .D(asr1_en_7_), .Q(asr2_rom_0__7_), .R(_225__bF_buf9), .S(1'b1) );
DFFSR DFFSR_137 ( .CLK(clk2_clkout_bF_buf22), .D(asr2_rom_6__0_), .Q(asr2_rom_7__0_), .R(_225__bF_buf8), .S(1'b1) );
DFFSR DFFSR_138 ( .CLK(clk2_clkout_bF_buf36), .D(asr2_rom_6__1_), .Q(asr2_rom_7__1_), .R(_225__bF_buf0), .S(1'b1) );
DFFSR DFFSR_139 ( .CLK(clk2_clkout_bF_buf25), .D(asr2_rom_6__2_), .Q(asr2_rom_7__2_), .R(_225__bF_buf1), .S(1'b1) );
DFFSR DFFSR_140 ( .CLK(clk2_clkout_bF_buf31), .D(asr2_rom_6__3_), .Q(asr2_rom_7__3_), .R(_225__bF_buf2), .S(1'b1) );
DFFSR DFFSR_141 ( .CLK(clk2_clkout_bF_buf3), .D(asr2_rom_6__4_), .Q(asr2_rom_7__4_), .R(_225__bF_buf0), .S(1'b1) );
DFFSR DFFSR_142 ( .CLK(clk2_clkout_bF_buf27), .D(asr2_rom_6__5_), .Q(asr2_rom_7__5_), .R(_225__bF_buf10), .S(1'b1) );
DFFSR DFFSR_143 ( .CLK(clk2_clkout_bF_buf22), .D(asr2_rom_6__6_), .Q(asr2_rom_7__6_), .R(_225__bF_buf8), .S(1'b1) );
DFFSR DFFSR_144 ( .CLK(clk2_clkout_bF_buf28), .D(asr2_rom_6__7_), .Q(asr2_rom_7__7_), .R(_225__bF_buf6), .S(1'b1) );
DFFSR DFFSR_145 ( .CLK(clk2_clkout_bF_buf17), .D(asr2_rom_1__0_), .Q(asr2_rom_2__0_), .R(_225__bF_buf3), .S(1'b1) );
DFFSR DFFSR_146 ( .CLK(clk2_clkout_bF_buf39), .D(asr2_rom_1__1_), .Q(asr2_rom_2__1_), .R(_225__bF_buf5), .S(1'b1) );
DFFSR DFFSR_147 ( .CLK(clk2_clkout_bF_buf25), .D(asr2_rom_1__2_), .Q(asr2_rom_2__2_), .R(_225__bF_buf1), .S(1'b1) );
DFFSR DFFSR_148 ( .CLK(clk2_clkout_bF_buf11), .D(asr2_rom_1__3_), .Q(asr2_rom_2__3_), .R(_225__bF_buf10), .S(1'b1) );
DFFSR DFFSR_149 ( .CLK(clk2_clkout_bF_buf32), .D(asr2_rom_1__4_), .Q(asr2_rom_2__4_), .R(_225__bF_buf8), .S(1'b1) );
DFFSR DFFSR_150 ( .CLK(clk2_clkout_bF_buf20), .D(asr2_rom_1__5_), .Q(asr2_rom_2__5_), .R(_225__bF_buf9), .S(1'b1) );
DFFSR DFFSR_151 ( .CLK(clk2_clkout_bF_buf28), .D(asr2_rom_1__6_), .Q(asr2_rom_2__6_), .R(_225__bF_buf6), .S(1'b1) );
DFFSR DFFSR_152 ( .CLK(clk2_clkout_bF_buf3), .D(asr2_rom_1__7_), .Q(asr2_rom_2__7_), .R(_225__bF_buf7), .S(1'b1) );
DFFSR DFFSR_153 ( .CLK(clk2_clkout_bF_buf40), .D(asr2_rom_0__0_), .Q(asr2_rom_1__0_), .R(_225__bF_buf3), .S(1'b1) );
DFFSR DFFSR_154 ( .CLK(clk2_clkout_bF_buf39), .D(asr2_rom_0__1_), .Q(asr2_rom_1__1_), .R(_225__bF_buf7), .S(1'b1) );
DFFSR DFFSR_155 ( .CLK(clk2_clkout_bF_buf20), .D(asr2_rom_0__2_), .Q(asr2_rom_1__2_), .R(_225__bF_buf9), .S(1'b1) );
DFFSR DFFSR_156 ( .CLK(clk2_clkout_bF_buf40), .D(asr2_rom_0__3_), .Q(asr2_rom_1__3_), .R(_225__bF_buf3), .S(1'b1) );
DFFSR DFFSR_157 ( .CLK(clk2_clkout_bF_buf28), .D(asr2_rom_0__4_), .Q(asr2_rom_1__4_), .R(_225__bF_buf4), .S(1'b1) );
DFFSR DFFSR_158 ( .CLK(clk2_clkout_bF_buf20), .D(asr2_rom_0__5_), .Q(asr2_rom_1__5_), .R(_225__bF_buf9), .S(1'b1) );
DFFSR DFFSR_159 ( .CLK(clk2_clkout_bF_buf22), .D(asr2_rom_0__6_), .Q(asr2_rom_1__6_), .R(_225__bF_buf1), .S(1'b1) );
DFFSR DFFSR_160 ( .CLK(clk2_clkout_bF_buf3), .D(asr2_rom_0__7_), .Q(asr2_rom_1__7_), .R(_225__bF_buf7), .S(1'b1) );
DFFSR DFFSR_161 ( .CLK(clk2_clkout_bF_buf40), .D(asr2_rom_2__0_), .Q(asr2_rom_3__0_), .R(_225__bF_buf3), .S(1'b1) );
DFFSR DFFSR_162 ( .CLK(clk2_clkout_bF_buf39), .D(asr2_rom_2__1_), .Q(asr2_rom_3__1_), .R(_225__bF_buf7), .S(1'b1) );
DFFSR DFFSR_163 ( .CLK(clk2_clkout_bF_buf13), .D(asr2_rom_2__2_), .Q(asr2_rom_3__2_), .R(_225__bF_buf4), .S(1'b1) );
DFFSR DFFSR_164 ( .CLK(clk2_clkout_bF_buf21), .D(asr2_rom_2__3_), .Q(asr2_rom_3__3_), .R(_225__bF_buf10), .S(1'b1) );
DFFSR DFFSR_165 ( .CLK(clk2_clkout_bF_buf32), .D(asr2_rom_2__4_), .Q(asr2_rom_3__4_), .R(_225__bF_buf8), .S(1'b1) );
DFFSR DFFSR_166 ( .CLK(clk2_clkout_bF_buf20), .D(asr2_rom_2__5_), .Q(asr2_rom_3__5_), .R(_225__bF_buf9), .S(1'b1) );
DFFSR DFFSR_167 ( .CLK(clk2_clkout_bF_buf32), .D(asr2_rom_2__6_), .Q(asr2_rom_3__6_), .R(_225__bF_buf6), .S(1'b1) );
DFFSR DFFSR_168 ( .CLK(clk2_clkout_bF_buf3), .D(asr2_rom_2__7_), .Q(asr2_rom_3__7_), .R(_225__bF_buf7), .S(1'b1) );
DFFSR DFFSR_169 ( .CLK(clk2_clkout_bF_buf31), .D(asr2_rom_3__0_), .Q(asr2_rom_4__0_), .R(_225__bF_buf1), .S(1'b1) );
DFFSR DFFSR_170 ( .CLK(clk2_clkout_bF_buf39), .D(asr2_rom_3__1_), .Q(asr2_rom_4__1_), .R(_225__bF_buf7), .S(1'b1) );
DFFSR DFFSR_171 ( .CLK(clk2_clkout_bF_buf13), .D(asr2_rom_3__2_), .Q(asr2_rom_4__2_), .R(_225__bF_buf9), .S(1'b1) );
DFFSR DFFSR_172 ( .CLK(clk2_clkout_bF_buf23), .D(asr2_rom_3__3_), .Q(asr2_rom_4__3_), .R(_225__bF_buf2), .S(1'b1) );
DFFSR DFFSR_173 ( .CLK(clk2_clkout_bF_buf28), .D(asr2_rom_3__4_), .Q(asr2_rom_4__4_), .R(_225__bF_buf6), .S(1'b1) );
DFFSR DFFSR_174 ( .CLK(clk2_clkout_bF_buf25), .D(asr2_rom_3__5_), .Q(asr2_rom_4__5_), .R(_225__bF_buf9), .S(1'b1) );
DFFSR DFFSR_175 ( .CLK(clk2_clkout_bF_buf32), .D(asr2_rom_3__6_), .Q(asr2_rom_4__6_), .R(_225__bF_buf6), .S(1'b1) );
DFFSR DFFSR_176 ( .CLK(clk2_clkout_bF_buf3), .D(asr2_rom_3__7_), .Q(asr2_rom_4__7_), .R(_225__bF_buf7), .S(1'b1) );
DFFSR DFFSR_177 ( .CLK(clk2_clkout_bF_buf22), .D(asr2_rom_5__0_), .Q(asr2_rom_6__0_), .R(_225__bF_buf1), .S(1'b1) );
DFFSR DFFSR_178 ( .CLK(clk2_clkout_bF_buf30), .D(asr2_rom_5__1_), .Q(asr2_rom_6__1_), .R(_225__bF_buf0), .S(1'b1) );
DFFSR DFFSR_179 ( .CLK(clk2_clkout_bF_buf20), .D(asr2_rom_5__2_), .Q(asr2_rom_6__2_), .R(_225__bF_buf9), .S(1'b1) );
DFFSR DFFSR_180 ( .CLK(clk2_clkout_bF_buf23), .D(asr2_rom_5__3_), .Q(asr2_rom_6__3_), .R(_225__bF_buf1), .S(1'b1) );
DFFSR DFFSR_181 ( .CLK(clk2_clkout_bF_buf30), .D(asr2_rom_5__4_), .Q(asr2_rom_6__4_), .R(_225__bF_buf0), .S(1'b1) );
DFFSR DFFSR_182 ( .CLK(clk2_clkout_bF_buf11), .D(asr2_rom_5__5_), .Q(asr2_rom_6__5_), .R(_225__bF_buf10), .S(1'b1) );
DFFSR DFFSR_183 ( .CLK(clk2_clkout_bF_buf8), .D(asr2_rom_5__6_), .Q(asr2_rom_6__6_), .R(_225__bF_buf8), .S(1'b1) );
DFFSR DFFSR_184 ( .CLK(clk2_clkout_bF_buf20), .D(asr2_rom_5__7_), .Q(asr2_rom_6__7_), .R(_225__bF_buf0), .S(1'b1) );
DFFSR DFFSR_185 ( .CLK(clk2_clkout_bF_buf25), .D(asr2_rom_4__0_), .Q(asr2_rom_5__0_), .R(_225__bF_buf1), .S(1'b1) );
DFFSR DFFSR_186 ( .CLK(clk2_clkout_bF_buf39), .D(asr2_rom_4__1_), .Q(asr2_rom_5__1_), .R(_225__bF_buf7), .S(1'b1) );
DFFSR DFFSR_187 ( .CLK(clk2_clkout_bF_buf13), .D(asr2_rom_4__2_), .Q(asr2_rom_5__2_), .R(_225__bF_buf4), .S(1'b1) );
DFFSR DFFSR_188 ( .CLK(clk2_clkout_bF_buf23), .D(asr2_rom_4__3_), .Q(asr2_rom_5__3_), .R(_225__bF_buf2), .S(1'b1) );
DFFSR DFFSR_189 ( .CLK(clk2_clkout_bF_buf30), .D(asr2_rom_4__4_), .Q(asr2_rom_5__4_), .R(_225__bF_buf0), .S(1'b1) );
DFFSR DFFSR_190 ( .CLK(clk2_clkout_bF_buf25), .D(asr2_rom_4__5_), .Q(asr2_rom_5__5_), .R(_225__bF_buf1), .S(1'b1) );
DFFSR DFFSR_191 ( .CLK(clk2_clkout_bF_buf32), .D(asr2_rom_4__6_), .Q(asr2_rom_5__6_), .R(_225__bF_buf6), .S(1'b1) );
DFFSR DFFSR_192 ( .CLK(clk2_clkout_bF_buf3), .D(asr2_rom_4__7_), .Q(asr2_rom_5__7_), .R(_225__bF_buf7), .S(1'b1) );
DFFSR DFFSR_193 ( .CLK(clk2_clkout_bF_buf8), .D(asr2_rom_7__0_), .Q(asr2_rom_8__0_), .R(_225__bF_buf8), .S(1'b1) );
DFFSR DFFSR_194 ( .CLK(clk2_clkout_bF_buf36), .D(asr2_rom_7__1_), .Q(asr2_rom_8__1_), .R(_225__bF_buf0), .S(1'b1) );
DFFSR DFFSR_195 ( .CLK(clk2_clkout_bF_buf31), .D(asr2_rom_7__2_), .Q(asr2_rom_8__2_), .R(_225__bF_buf1), .S(1'b1) );
DFFSR DFFSR_196 ( .CLK(clk2_clkout_bF_buf21), .D(asr2_rom_7__3_), .Q(asr2_rom_8__3_), .R(_225__bF_buf2), .S(1'b1) );
DFFSR DFFSR_197 ( .CLK(clk2_clkout_bF_buf2), .D(asr2_rom_7__4_), .Q(asr2_rom_8__4_), .R(_225__bF_buf7), .S(1'b1) );
DFFSR DFFSR_198 ( .CLK(clk2_clkout_bF_buf21), .D(asr2_rom_7__5_), .Q(asr2_rom_8__5_), .R(_225__bF_buf2), .S(1'b1) );
DFFSR DFFSR_199 ( .CLK(clk2_clkout_bF_buf22), .D(asr2_rom_7__6_), .Q(asr2_rom_8__6_), .R(_225__bF_buf4), .S(1'b1) );
DFFSR DFFSR_200 ( .CLK(clk2_clkout_bF_buf28), .D(asr2_rom_7__7_), .Q(asr2_rom_8__7_), .R(_225__bF_buf6), .S(1'b1) );
DFFSR DFFSR_201 ( .CLK(clk2_clkout_bF_buf8), .D(asr2_rom_8__0_), .Q(asr2_rom_9__0_), .R(_225__bF_buf8), .S(1'b1) );
DFFSR DFFSR_202 ( .CLK(clk2_clkout_bF_buf30), .D(asr2_rom_8__1_), .Q(asr2_rom_9__1_), .R(_225__bF_buf0), .S(1'b1) );
DFFSR DFFSR_203 ( .CLK(clk2_clkout_bF_buf23), .D(asr2_rom_8__2_), .Q(asr2_rom_9__2_), .R(_225__bF_buf2), .S(1'b1) );
DFFSR DFFSR_204 ( .CLK(clk2_clkout_bF_buf27), .D(asr2_rom_8__3_), .Q(asr2_rom_9__3_), .R(_225__bF_buf10), .S(1'b1) );
DFFSR DFFSR_205 ( .CLK(clk2_clkout_bF_buf20), .D(asr2_rom_8__4_), .Q(asr2_rom_9__4_), .R(_225__bF_buf9), .S(1'b1) );
DFFSR DFFSR_206 ( .CLK(clk2_clkout_bF_buf21), .D(asr2_rom_8__5_), .Q(asr2_rom_9__5_), .R(_225__bF_buf10), .S(1'b1) );
DFFSR DFFSR_207 ( .CLK(clk2_clkout_bF_buf22), .D(asr2_rom_8__6_), .Q(asr2_rom_9__6_), .R(_225__bF_buf4), .S(1'b1) );
DFFSR DFFSR_208 ( .CLK(clk2_clkout_bF_buf28), .D(asr2_rom_8__7_), .Q(asr2_rom_9__7_), .R(_225__bF_buf6), .S(1'b1) );
DFFSR DFFSR_209 ( .CLK(clk2_clkout_bF_buf8), .D(asr2_rom_9__0_), .Q(asr2_rom_10__0_), .R(_225__bF_buf8), .S(1'b1) );
DFFSR DFFSR_210 ( .CLK(clk2_clkout_bF_buf41), .D(asr2_rom_9__1_), .Q(asr2_rom_10__1_), .R(_225__bF_buf5), .S(1'b1) );
DFFSR DFFSR_211 ( .CLK(clk2_clkout_bF_buf31), .D(asr2_rom_9__2_), .Q(asr2_rom_10__2_), .R(_225__bF_buf2), .S(1'b1) );
DFFSR DFFSR_212 ( .CLK(clk2_clkout_bF_buf11), .D(asr2_rom_9__3_), .Q(asr2_rom_10__3_), .R(_225__bF_buf10), .S(1'b1) );
DFFSR DFFSR_213 ( .CLK(clk2_clkout_bF_buf30), .D(asr2_rom_9__4_), .Q(asr2_rom_10__4_), .R(_225__bF_buf0), .S(1'b1) );
DFFSR DFFSR_214 ( .CLK(clk2_clkout_bF_buf17), .D(asr2_rom_9__5_), .Q(asr2_rom_10__5_), .R(_225__bF_buf10), .S(1'b1) );
DFFSR DFFSR_215 ( .CLK(clk2_clkout_bF_buf13), .D(asr2_rom_9__6_), .Q(asr2_rom_10__6_), .R(_225__bF_buf4), .S(1'b1) );
DFFSR DFFSR_216 ( .CLK(clk2_clkout_bF_buf32), .D(asr2_rom_9__7_), .Q(asr2_rom_10__7_), .R(_225__bF_buf6), .S(1'b1) );
DFFSR DFFSR_217 ( .CLK(clk2_clkout_bF_buf8), .D(asr2_rom_10__0_), .Q(asr2_rom_11__0_), .R(_225__bF_buf8), .S(1'b1) );
DFFSR DFFSR_218 ( .CLK(clk2_clkout_bF_buf41), .D(asr2_rom_10__1_), .Q(asr2_rom_11__1_), .R(_225__bF_buf5), .S(1'b1) );
DFFSR DFFSR_219 ( .CLK(clk2_clkout_bF_buf17), .D(asr2_rom_10__2_), .Q(asr2_rom_11__2_), .R(_225__bF_buf10), .S(1'b1) );
DFFSR DFFSR_220 ( .CLK(clk2_clkout_bF_buf11), .D(asr2_rom_10__3_), .Q(asr2_rom_11__3_), .R(_225__bF_buf10), .S(1'b1) );
DFFSR DFFSR_221 ( .CLK(clk2_clkout_bF_buf30), .D(asr2_rom_10__4_), .Q(asr2_rom_11__4_), .R(_225__bF_buf0), .S(1'b1) );
DFFSR DFFSR_222 ( .CLK(clk2_clkout_bF_buf17), .D(asr2_rom_10__5_), .Q(asr2_rom_11__5_), .R(_225__bF_buf10), .S(1'b1) );
DFFSR DFFSR_223 ( .CLK(clk2_clkout_bF_buf13), .D(asr2_rom_10__6_), .Q(asr2_rom_11__6_), .R(_225__bF_buf4), .S(1'b1) );
DFFSR DFFSR_224 ( .CLK(clk2_clkout_bF_buf32), .D(asr2_rom_10__7_), .Q(asr2_rom_11__7_), .R(_225__bF_buf6), .S(1'b1) );
DFFSR DFFSR_225 ( .CLK(clk2_clkout_bF_buf8), .D(asr2_rom_11__0_), .Q(asr2_rom_12__0_), .R(_225__bF_buf8), .S(1'b1) );
DFFSR DFFSR_226 ( .CLK(clk2_clkout_bF_buf12), .D(asr2_rom_11__1_), .Q(asr2_rom_12__1_), .R(_225__bF_buf5), .S(1'b1) );
DFFSR DFFSR_227 ( .CLK(clk2_clkout_bF_buf21), .D(asr2_rom_11__2_), .Q(asr2_rom_12__2_), .R(_225__bF_buf2), .S(1'b1) );
DFFSR DFFSR_228 ( .CLK(clk2_clkout_bF_buf21), .D(asr2_rom_11__3_), .Q(asr2_rom_12__3_), .R(_225__bF_buf2), .S(1'b1) );
DFFSR DFFSR_229 ( .CLK(clk2_clkout_bF_buf30), .D(asr2_rom_11__4_), .Q(asr2_rom_12__4_), .R(_225__bF_buf0), .S(1'b1) );
DFFSR DFFSR_230 ( .CLK(clk2_clkout_bF_buf17), .D(asr2_rom_11__5_), .Q(asr2_rom_12__5_), .R(_225__bF_buf10), .S(1'b1) );
DFFSR DFFSR_231 ( .CLK(clk2_clkout_bF_buf13), .D(asr2_rom_11__6_), .Q(asr2_rom_12__6_), .R(_225__bF_buf4), .S(1'b1) );
DFFSR DFFSR_232 ( .CLK(clk2_clkout_bF_buf28), .D(asr2_rom_11__7_), .Q(asr2_rom_12__7_), .R(_225__bF_buf6), .S(1'b1) );
DFFSR DFFSR_233 ( .CLK(clk2_clkout_bF_buf40), .D(asr2_rom_12__0_), .Q(asr2_rom_13__0_), .R(_225__bF_buf8), .S(1'b1) );
DFFSR DFFSR_234 ( .CLK(clk2_clkout_bF_buf12), .D(asr2_rom_12__1_), .Q(asr2_rom_13__1_), .R(_225__bF_buf5), .S(1'b1) );
DFFSR DFFSR_235 ( .CLK(clk2_clkout_bF_buf40), .D(asr2_rom_12__2_), .Q(asr2_rom_13__2_), .R(_225__bF_buf3), .S(1'b1) );
DFFSR DFFSR_236 ( .CLK(clk2_clkout_bF_buf21), .D(asr2_rom_12__3_), .Q(asr2_rom_13__3_), .R(_225__bF_buf2), .S(1'b1) );
DFFSR DFFSR_237 ( .CLK(clk2_clkout_bF_buf36), .D(asr2_rom_12__4_), .Q(asr2_rom_13__4_), .R(_225__bF_buf4), .S(1'b1) );
DFFSR DFFSR_238 ( .CLK(clk2_clkout_bF_buf17), .D(asr2_rom_12__5_), .Q(asr2_rom_13__5_), .R(_225__bF_buf3), .S(1'b1) );
DFFSR DFFSR_239 ( .CLK(clk2_clkout_bF_buf36), .D(asr2_rom_12__6_), .Q(asr2_rom_13__6_), .R(_225__bF_buf6), .S(1'b1) );
DFFSR DFFSR_240 ( .CLK(clk2_clkout_bF_buf36), .D(asr2_rom_12__7_), .Q(asr2_rom_13__7_), .R(_225__bF_buf4), .S(1'b1) );
DFFSR DFFSR_241 ( .CLK(clk2_clkout_bF_buf40), .D(asr2_rom_13__0_), .Q(asr2_rom_14__0_), .R(_225__bF_buf3), .S(1'b1) );
DFFSR DFFSR_242 ( .CLK(clk2_clkout_bF_buf12), .D(asr2_rom_13__1_), .Q(asr2_rom_14__1_), .R(_225__bF_buf5), .S(1'b1) );
DFFSR DFFSR_243 ( .CLK(clk2_clkout_bF_buf31), .D(asr2_rom_13__2_), .Q(asr2_rom_14__2_), .R(_225__bF_buf3), .S(1'b1) );
DFFSR DFFSR_244 ( .CLK(clk2_clkout_bF_buf25), .D(asr2_rom_13__3_), .Q(asr2_rom_14__3_), .R(_225__bF_buf1), .S(1'b1) );
DFFSR DFFSR_245 ( .CLK(clk2_clkout_bF_buf36), .D(asr2_rom_13__4_), .Q(asr2_rom_14__4_), .R(_225__bF_buf4), .S(1'b1) );
DFFSR DFFSR_246 ( .CLK(clk2_clkout_bF_buf31), .D(asr2_rom_13__5_), .Q(asr2_rom_14__5_), .R(_225__bF_buf3), .S(1'b1) );
DFFSR DFFSR_247 ( .CLK(clk2_clkout_bF_buf39), .D(asr2_rom_13__6_), .Q(asr2_rom_14__6_), .R(_225__bF_buf5), .S(1'b1) );
DFFSR DFFSR_248 ( .CLK(clk2_clkout_bF_buf41), .D(asr2_rom_13__7_), .Q(asr2_rom_14__7_), .R(_225__bF_buf5), .S(1'b1) );
DFFSR DFFSR_249 ( .CLK(clk2_clkout_bF_buf40), .D(asr2_rom_14__0_), .Q(asr2_en_0_), .R(_225__bF_buf3), .S(1'b1) );
DFFSR DFFSR_250 ( .CLK(clk2_clkout_bF_buf19), .D(asr2_rom_14__1_), .Q(asr2_en_1_), .R(_225__bF_buf5), .S(1'b1) );
DFFSR DFFSR_251 ( .CLK(clk2_clkout_bF_buf22), .D(asr2_rom_14__2_), .Q(asr2_en_2_), .R(_225__bF_buf8), .S(1'b1) );
DFFSR DFFSR_252 ( .CLK(clk2_clkout_bF_buf24), .D(asr2_rom_14__3_), .Q(asr2_en_3_), .R(_225__bF_buf9), .S(1'b1) );
DFFSR DFFSR_253 ( .CLK(clk2_clkout_bF_buf36), .D(asr2_rom_14__4_), .Q(asr2_en_4_), .R(_225__bF_buf4), .S(1'b1) );
DFFSR DFFSR_254 ( .CLK(clk2_clkout_bF_buf25), .D(asr2_rom_14__5_), .Q(asr2_en_5_), .R(_225__bF_buf1), .S(1'b1) );
DFFSR DFFSR_255 ( .CLK(clk2_clkout_bF_buf41), .D(asr2_rom_14__6_), .Q(asr2_en_6_), .R(_225__bF_buf5), .S(1'b1) );
DFFSR DFFSR_256 ( .CLK(clk2_clkout_bF_buf19), .D(asr2_rom_14__7_), .Q(asr2_en_7_), .R(_225__bF_buf5), .S(1'b1) );
NOR2X1 NOR2X1_59 ( .A(rst_bF_buf2), .B(clk2_div_0_), .Y(_451__0_) );
INVX1 INVX1_119 ( .A(rst_bF_buf1), .Y(_452_) );
OAI21X1 OAI21X1_17 ( .A(clk2_div_0_), .B(clk2_div_1_), .C(_452_), .Y(_453_) );
AOI21X1 AOI21X1_1 ( .A(clk2_div_0_), .B(clk2_div_1_), .C(_453_), .Y(_451__1_) );
NAND3X1 NAND3X1_129 ( .A(clk2_div_0_), .B(clk2_div_1_), .C(clk2_div_2_), .Y(_454_) );
INVX1 INVX1_120 ( .A(clk2_div_2_), .Y(_455_) );
NAND2X1 NAND2X1_53 ( .A(clk2_div_0_), .B(clk2_div_1_), .Y(_456_) );
AOI21X1 AOI21X1_2 ( .A(_456_), .B(_455_), .C(rst_bF_buf1), .Y(_457_) );
AND2X2 AND2X2_27 ( .A(_457_), .B(_454_), .Y(_451__2_) );
AOI21X1 AOI21X1_3 ( .A(_454_), .B(clk2_clkout_bF_buf10), .C(rst_bF_buf2), .Y(_458_) );
OAI21X1 OAI21X1_18 ( .A(clk2_clkout_bF_buf10), .B(_454_), .C(_458_), .Y(_450_) );
DFFPOSX1 DFFPOSX1_1 ( .CLK(clk_bF_buf0), .D(_450_), .Q(clk2_clkout) );
DFFPOSX1 DFFPOSX1_2 ( .CLK(clk_bF_buf0), .D(_451__0_), .Q(clk2_div_0_) );
DFFPOSX1 DFFPOSX1_3 ( .CLK(clk_bF_buf0), .D(_451__1_), .Q(clk2_div_1_) );
DFFPOSX1 DFFPOSX1_4 ( .CLK(clk_bF_buf5), .D(_451__2_), .Q(clk2_div_2_) );
OR2X2 OR2X2_1 ( .A(counterup_counter_1_), .B(counterup_counter_0_bF_buf0_), .Y(_462_) );
INVX1 INVX1_121 ( .A(counterup_counter_3_), .Y(_463_) );
INVX1 INVX1_122 ( .A(counterup_counter_2_), .Y(_464_) );
INVX1 INVX1_123 ( .A(rst_bF_buf2), .Y(_460_) );
NAND3X1 NAND3X1_130 ( .A(_463_), .B(_464_), .C(_460_), .Y(_461_) );
NOR2X1 NOR2X1_60 ( .A(_462_), .B(_461_), .Y(_459_) );
DFFPOSX1 DFFPOSX1_5 ( .CLK(clk_bF_buf5), .D(_459_), .Q(comp_dataout) );
INVX1 INVX1_124 ( .A(rst_bF_buf2), .Y(_466_) );
NAND2X1 NAND2X1_54 ( .A(counterdown_counter_0_), .B(_466_), .Y(_465__0_) );
AOI21X1 AOI21X1_4 ( .A(counterdown_counter_0_), .B(counterdown_counter_1_), .C(rst_bF_buf0), .Y(_467_) );
OAI21X1 OAI21X1_19 ( .A(counterdown_counter_0_), .B(counterdown_counter_1_), .C(_467_), .Y(_465__1_) );
INVX1 INVX1_125 ( .A(counterdown_counter_0_), .Y(_468_) );
INVX1 INVX1_126 ( .A(counterdown_counter_1_), .Y(_469_) );
INVX1 INVX1_127 ( .A(counterdown_counter_2_), .Y(_470_) );
NAND3X1 NAND3X1_131 ( .A(_468_), .B(_469_), .C(_470_), .Y(_471_) );
OAI21X1 OAI21X1_20 ( .A(counterdown_counter_0_), .B(counterdown_counter_1_), .C(counterdown_counter_2_), .Y(_472_) );
NAND3X1 NAND3X1_132 ( .A(_466_), .B(_472_), .C(_471_), .Y(_465__2_) );
NAND2X1 NAND2X1_55 ( .A(counterdown_counter_3_), .B(_471_), .Y(_473_) );
INVX1 INVX1_128 ( .A(counterdown_counter_3_), .Y(_474_) );
NOR2X1 NOR2X1_61 ( .A(counterdown_counter_0_), .B(counterdown_counter_1_), .Y(_475_) );
NAND3X1 NAND3X1_133 ( .A(_470_), .B(_474_), .C(_475_), .Y(_476_) );
NAND3X1 NAND3X1_134 ( .A(_466_), .B(_476_), .C(_473_), .Y(_465__3_) );
DFFPOSX1 DFFPOSX1_6 ( .CLK(clk_bF_buf6), .D(_465__0_), .Q(counterdown_counter_0_) );
DFFPOSX1 DFFPOSX1_7 ( .CLK(clk_bF_buf3), .D(_465__1_), .Q(counterdown_counter_1_) );
DFFPOSX1 DFFPOSX1_8 ( .CLK(clk_bF_buf3), .D(_465__2_), .Q(counterdown_counter_2_) );
DFFPOSX1 DFFPOSX1_9 ( .CLK(clk_bF_buf6), .D(_465__3_), .Q(counterdown_counter_3_) );
NOR2X1 NOR2X1_62 ( .A(counterup_counter_0_bF_buf3_), .B(rst_bF_buf4), .Y(_477__0_) );
AND2X2 AND2X2_28 ( .A(counterup_counter_0_bF_buf2_), .B(counterup_counter_1_), .Y(_478_) );
INVX1 INVX1_129 ( .A(rst_bF_buf5), .Y(_479_) );
OAI21X1 OAI21X1_21 ( .A(counterup_counter_0_bF_buf1_), .B(counterup_counter_1_), .C(_479_), .Y(_480_) );
NOR2X1 NOR2X1_63 ( .A(_478_), .B(_480_), .Y(_477__1_) );
AOI21X1 AOI21X1_5 ( .A(counterup_counter_0_bF_buf0_), .B(counterup_counter_1_), .C(counterup_counter_2_), .Y(_481_) );
NAND3X1 NAND3X1_135 ( .A(counterup_counter_0_bF_buf3_), .B(counterup_counter_1_), .C(counterup_counter_2_), .Y(_482_) );
NAND2X1 NAND2X1_56 ( .A(_479_), .B(_482_), .Y(_483_) );
NOR2X1 NOR2X1_64 ( .A(_481_), .B(_483_), .Y(_477__2_) );
NAND2X1 NAND2X1_57 ( .A(counterup_counter_3_), .B(_482_), .Y(_484_) );
INVX1 INVX1_130 ( .A(counterup_counter_3_), .Y(_485_) );
NAND3X1 NAND3X1_136 ( .A(counterup_counter_2_), .B(_485_), .C(_478_), .Y(_486_) );
AOI21X1 AOI21X1_6 ( .A(_486_), .B(_484_), .C(rst_bF_buf2), .Y(_477__3_) );
DFFPOSX1 DFFPOSX1_10 ( .CLK(clk_bF_buf6), .D(_477__0_), .Q(counterup_counter_0_) );
DFFPOSX1 DFFPOSX1_11 ( .CLK(clk_bF_buf3), .D(_477__1_), .Q(counterup_counter_1_) );
DFFPOSX1 DFFPOSX1_12 ( .CLK(clk_bF_buf1), .D(_477__2_), .Q(counterup_counter_2_) );
DFFPOSX1 DFFPOSX1_13 ( .CLK(clk_bF_buf6), .D(_477__3_), .Q(counterup_counter_3_) );
NAND2X1 NAND2X1_58 ( .A(rom1_data_0_bF_buf3_), .B(sumador_res_0_), .Y(_734_) );
INVX1 INVX1_131 ( .A(mac1_reset_bF_buf3), .Y(_745_) );
NAND2X1 NAND2X1_59 ( .A(mac1_dataout_0_), .B(_745_), .Y(_756_) );
XOR2X1 XOR2X1_1 ( .A(_756_), .B(_734_), .Y(_487__0_) );
INVX1 INVX1_132 ( .A(rom1_data_0_bF_buf2_), .Y(_777_) );
INVX1 INVX1_133 ( .A(sumador_res_0_), .Y(_788_) );
INVX1 INVX1_134 ( .A(sumador_res_1_), .Y(_795_) );
INVX1 INVX1_135 ( .A(rom1_data_1_), .Y(_796_) );
OAI22X1 OAI22X1_49 ( .A(_777_), .B(_795_), .C(_788_), .D(_796_), .Y(_797_) );
NAND2X1 NAND2X1_60 ( .A(sumador_res_1_), .B(rom1_data_1_), .Y(_798_) );
OAI21X1 OAI21X1_22 ( .A(_734_), .B(_798_), .C(_797_), .Y(_799_) );
NAND3X1 NAND3X1_137 ( .A(rom1_data_0_bF_buf1_), .B(sumador_res_0_), .C(mac1_dataout_0_), .Y(_800_) );
INVX1 INVX1_136 ( .A(_800_), .Y(_801_) );
INVX1 INVX1_137 ( .A(mac1_dataout_1_), .Y(_802_) );
XOR2X1 XOR2X1_2 ( .A(_799_), .B(_802_), .Y(_803_) );
NAND2X1 NAND2X1_61 ( .A(_801_), .B(_803_), .Y(_804_) );
OR2X2 OR2X2_2 ( .A(_803_), .B(_801_), .Y(_805_) );
NAND3X1 NAND3X1_138 ( .A(_745_), .B(_804_), .C(_805_), .Y(_806_) );
OAI21X1 OAI21X1_23 ( .A(_745_), .B(_799_), .C(_806_), .Y(_487__1_) );
NAND2X1 NAND2X1_62 ( .A(sumador_res_0_), .B(rom1_data_2_), .Y(_807_) );
INVX1 INVX1_138 ( .A(_807_), .Y(_808_) );
AND2X2 AND2X2_29 ( .A(rom1_data_0_bF_buf0_), .B(sumador_res_2_), .Y(_809_) );
NAND3X1 NAND3X1_139 ( .A(sumador_res_1_), .B(rom1_data_1_), .C(_809_), .Y(_810_) );
AOI22X1 AOI22X1_17 ( .A(rom1_data_0_bF_buf3_), .B(sumador_res_2_), .C(sumador_res_1_), .D(rom1_data_1_), .Y(_811_) );
INVX1 INVX1_139 ( .A(_811_), .Y(_812_) );
NAND3X1 NAND3X1_140 ( .A(_812_), .B(_808_), .C(_810_), .Y(_813_) );
NAND2X1 NAND2X1_63 ( .A(rom1_data_0_bF_buf2_), .B(sumador_res_2_), .Y(_814_) );
NOR2X1 NOR2X1_65 ( .A(_798_), .B(_814_), .Y(_815_) );
OAI21X1 OAI21X1_24 ( .A(_811_), .B(_815_), .C(_807_), .Y(_816_) );
NAND2X1 NAND2X1_64 ( .A(_813_), .B(_816_), .Y(_817_) );
OAI21X1 OAI21X1_25 ( .A(_734_), .B(_798_), .C(_817_), .Y(_818_) );
NOR2X1 NOR2X1_66 ( .A(_734_), .B(_798_), .Y(_819_) );
NAND3X1 NAND3X1_141 ( .A(_819_), .B(_813_), .C(_816_), .Y(_820_) );
NAND2X1 NAND2X1_65 ( .A(_820_), .B(_818_), .Y(_821_) );
OAI21X1 OAI21X1_26 ( .A(_802_), .B(_799_), .C(_804_), .Y(_822_) );
INVX1 INVX1_140 ( .A(_822_), .Y(_823_) );
NAND3X1 NAND3X1_142 ( .A(mac1_dataout_2_), .B(_820_), .C(_818_), .Y(_824_) );
INVX1 INVX1_141 ( .A(_824_), .Y(_825_) );
AOI21X1 AOI21X1_7 ( .A(_818_), .B(_820_), .C(mac1_dataout_2_), .Y(_826_) );
NOR2X1 NOR2X1_67 ( .A(_826_), .B(_825_), .Y(_827_) );
AND2X2 AND2X2_30 ( .A(_827_), .B(_823_), .Y(_828_) );
NOR2X1 NOR2X1_68 ( .A(_823_), .B(_827_), .Y(_829_) );
OAI21X1 OAI21X1_27 ( .A(_829_), .B(_828_), .C(_745_), .Y(_830_) );
OAI21X1 OAI21X1_28 ( .A(_745_), .B(_821_), .C(_830_), .Y(_487__2_) );
OAI21X1 OAI21X1_29 ( .A(_826_), .B(_823_), .C(_824_), .Y(_831_) );
INVX1 INVX1_142 ( .A(_820_), .Y(_832_) );
NAND2X1 NAND2X1_66 ( .A(sumador_res_0_), .B(rom1_data_3_), .Y(_833_) );
INVX1 INVX1_143 ( .A(_833_), .Y(_834_) );
OAI21X1 OAI21X1_30 ( .A(_807_), .B(_811_), .C(_810_), .Y(_835_) );
NAND2X1 NAND2X1_67 ( .A(sumador_res_1_), .B(rom1_data_2_), .Y(_836_) );
INVX1 INVX1_144 ( .A(_836_), .Y(_837_) );
AND2X2 AND2X2_31 ( .A(rom1_data_1_), .B(sumador_res_2_), .Y(_838_) );
AND2X2 AND2X2_32 ( .A(rom1_data_0_bF_buf1_), .B(sumador_res_3_), .Y(_839_) );
NAND2X1 NAND2X1_68 ( .A(_838_), .B(_839_), .Y(_840_) );
INVX1 INVX1_145 ( .A(sumador_res_2_), .Y(_841_) );
NAND2X1 NAND2X1_69 ( .A(rom1_data_0_bF_buf0_), .B(sumador_res_3_), .Y(_842_) );
OAI21X1 OAI21X1_31 ( .A(_796_), .B(_841_), .C(_842_), .Y(_843_) );
NAND3X1 NAND3X1_143 ( .A(_843_), .B(_837_), .C(_840_), .Y(_844_) );
OAI21X1 OAI21X1_32 ( .A(_796_), .B(_841_), .C(_839_), .Y(_845_) );
INVX1 INVX1_146 ( .A(sumador_res_3_), .Y(_846_) );
OAI21X1 OAI21X1_33 ( .A(_777_), .B(_846_), .C(_838_), .Y(_847_) );
NAND3X1 NAND3X1_144 ( .A(_836_), .B(_845_), .C(_847_), .Y(_848_) );
NAND3X1 NAND3X1_145 ( .A(_844_), .B(_835_), .C(_848_), .Y(_849_) );
AOI21X1 AOI21X1_8 ( .A(_808_), .B(_812_), .C(_815_), .Y(_850_) );
NAND3X1 NAND3X1_146 ( .A(_836_), .B(_843_), .C(_840_), .Y(_851_) );
NAND3X1 NAND3X1_147 ( .A(_837_), .B(_845_), .C(_847_), .Y(_852_) );
NAND3X1 NAND3X1_148 ( .A(_851_), .B(_852_), .C(_850_), .Y(_488_) );
NAND3X1 NAND3X1_149 ( .A(_834_), .B(_849_), .C(_488_), .Y(_489_) );
NAND3X1 NAND3X1_150 ( .A(_844_), .B(_848_), .C(_850_), .Y(_490_) );
NAND3X1 NAND3X1_151 ( .A(_851_), .B(_835_), .C(_852_), .Y(_491_) );
NAND3X1 NAND3X1_152 ( .A(_833_), .B(_491_), .C(_490_), .Y(_492_) );
AOI21X1 AOI21X1_9 ( .A(_489_), .B(_492_), .C(_832_), .Y(_493_) );
INVX1 INVX1_147 ( .A(_493_), .Y(_494_) );
NAND3X1 NAND3X1_153 ( .A(_832_), .B(_489_), .C(_492_), .Y(_495_) );
NAND3X1 NAND3X1_154 ( .A(mac1_dataout_3_), .B(_495_), .C(_494_), .Y(_496_) );
INVX1 INVX1_148 ( .A(mac1_dataout_3_), .Y(_497_) );
INVX1 INVX1_149 ( .A(_495_), .Y(_498_) );
OAI21X1 OAI21X1_34 ( .A(_493_), .B(_498_), .C(_497_), .Y(_499_) );
NAND2X1 NAND2X1_70 ( .A(_496_), .B(_499_), .Y(_500_) );
XOR2X1 XOR2X1_3 ( .A(_500_), .B(_831_), .Y(_501_) );
NAND3X1 NAND3X1_155 ( .A(mac1_reset_bF_buf1), .B(_495_), .C(_494_), .Y(_502_) );
OAI21X1 OAI21X1_35 ( .A(mac1_reset_bF_buf2), .B(_501_), .C(_502_), .Y(_487__3_) );
NAND2X1 NAND2X1_71 ( .A(sumador_res_1_), .B(rom1_data_4_), .Y(_503_) );
INVX1 INVX1_150 ( .A(rom1_data_4_), .Y(_504_) );
NAND2X1 NAND2X1_72 ( .A(sumador_res_1_), .B(rom1_data_3_), .Y(_505_) );
OAI21X1 OAI21X1_36 ( .A(_788_), .B(_504_), .C(_505_), .Y(_506_) );
OAI21X1 OAI21X1_37 ( .A(_833_), .B(_503_), .C(_506_), .Y(_507_) );
AOI22X1 AOI22X1_18 ( .A(rom1_data_0_bF_buf3_), .B(sumador_res_3_), .C(rom1_data_1_), .D(sumador_res_2_), .Y(_508_) );
OAI21X1 OAI21X1_38 ( .A(_836_), .B(_508_), .C(_840_), .Y(_509_) );
NAND2X1 NAND2X1_73 ( .A(sumador_res_2_), .B(rom1_data_2_), .Y(_510_) );
INVX1 INVX1_151 ( .A(_510_), .Y(_511_) );
AND2X2 AND2X2_33 ( .A(rom1_data_1_), .B(sumador_res_4_), .Y(_512_) );
NAND2X1 NAND2X1_74 ( .A(_839_), .B(_512_), .Y(_513_) );
NAND2X1 NAND2X1_75 ( .A(rom1_data_1_), .B(sumador_res_3_), .Y(_514_) );
NAND2X1 NAND2X1_76 ( .A(rom1_data_0_bF_buf2_), .B(sumador_res_4_), .Y(_515_) );
NAND2X1 NAND2X1_77 ( .A(_514_), .B(_515_), .Y(_516_) );
NAND3X1 NAND3X1_156 ( .A(_511_), .B(_516_), .C(_513_), .Y(_517_) );
NAND3X1 NAND3X1_157 ( .A(rom1_data_0_bF_buf1_), .B(sumador_res_4_), .C(_514_), .Y(_518_) );
AND2X2 AND2X2_34 ( .A(rom1_data_1_), .B(sumador_res_3_), .Y(_519_) );
NAND2X1 NAND2X1_78 ( .A(_515_), .B(_519_), .Y(_520_) );
NAND3X1 NAND3X1_158 ( .A(_510_), .B(_518_), .C(_520_), .Y(_521_) );
NAND3X1 NAND3X1_159 ( .A(_509_), .B(_517_), .C(_521_), .Y(_522_) );
AOI22X1 AOI22X1_19 ( .A(_809_), .B(_519_), .C(_843_), .D(_837_), .Y(_523_) );
NAND3X1 NAND3X1_160 ( .A(_510_), .B(_516_), .C(_513_), .Y(_524_) );
NAND3X1 NAND3X1_161 ( .A(_511_), .B(_518_), .C(_520_), .Y(_525_) );
NAND3X1 NAND3X1_162 ( .A(_525_), .B(_524_), .C(_523_), .Y(_526_) );
NAND3X1 NAND3X1_163 ( .A(_507_), .B(_522_), .C(_526_), .Y(_527_) );
INVX1 INVX1_152 ( .A(_507_), .Y(_528_) );
AOI21X1 AOI21X1_10 ( .A(_524_), .B(_525_), .C(_523_), .Y(_529_) );
AOI21X1 AOI21X1_11 ( .A(_517_), .B(_521_), .C(_509_), .Y(_530_) );
OAI21X1 OAI21X1_39 ( .A(_530_), .B(_529_), .C(_528_), .Y(_531_) );
AOI22X1 AOI22X1_20 ( .A(_849_), .B(_489_), .C(_531_), .D(_527_), .Y(_532_) );
AOI21X1 AOI21X1_12 ( .A(_848_), .B(_844_), .C(_835_), .Y(_533_) );
OAI21X1 OAI21X1_40 ( .A(_833_), .B(_533_), .C(_849_), .Y(_534_) );
NAND3X1 NAND3X1_164 ( .A(_528_), .B(_522_), .C(_526_), .Y(_535_) );
OAI21X1 OAI21X1_41 ( .A(_530_), .B(_529_), .C(_507_), .Y(_536_) );
AOI21X1 AOI21X1_13 ( .A(_535_), .B(_536_), .C(_534_), .Y(_537_) );
OAI21X1 OAI21X1_42 ( .A(_532_), .B(_537_), .C(_495_), .Y(_538_) );
NAND3X1 NAND3X1_165 ( .A(_535_), .B(_536_), .C(_534_), .Y(_539_) );
AOI21X1 AOI21X1_14 ( .A(_851_), .B(_852_), .C(_850_), .Y(_540_) );
AOI21X1 AOI21X1_15 ( .A(_834_), .B(_488_), .C(_540_), .Y(_541_) );
NAND3X1 NAND3X1_166 ( .A(_527_), .B(_531_), .C(_541_), .Y(_542_) );
NAND3X1 NAND3X1_167 ( .A(_539_), .B(_542_), .C(_498_), .Y(_543_) );
NAND2X1 NAND2X1_79 ( .A(_538_), .B(_543_), .Y(_544_) );
INVX1 INVX1_153 ( .A(_826_), .Y(_545_) );
AOI21X1 AOI21X1_16 ( .A(_545_), .B(_822_), .C(_825_), .Y(_546_) );
AOI21X1 AOI21X1_17 ( .A(_494_), .B(_495_), .C(mac1_dataout_3_), .Y(_547_) );
OAI21X1 OAI21X1_43 ( .A(_546_), .B(_547_), .C(_496_), .Y(_548_) );
NAND3X1 NAND3X1_168 ( .A(mac1_dataout_4_), .B(_538_), .C(_543_), .Y(_549_) );
INVX1 INVX1_154 ( .A(mac1_dataout_4_), .Y(_550_) );
NAND2X1 NAND2X1_80 ( .A(_550_), .B(_544_), .Y(_551_) );
NAND3X1 NAND3X1_169 ( .A(_549_), .B(_548_), .C(_551_), .Y(_552_) );
INVX1 INVX1_155 ( .A(_496_), .Y(_553_) );
AOI21X1 AOI21X1_18 ( .A(_499_), .B(_831_), .C(_553_), .Y(_554_) );
INVX1 INVX1_156 ( .A(_549_), .Y(_555_) );
AOI21X1 AOI21X1_19 ( .A(_543_), .B(_538_), .C(mac1_dataout_4_), .Y(_556_) );
OAI21X1 OAI21X1_44 ( .A(_556_), .B(_555_), .C(_554_), .Y(_557_) );
NAND3X1 NAND3X1_170 ( .A(_745_), .B(_552_), .C(_557_), .Y(_558_) );
OAI21X1 OAI21X1_45 ( .A(_745_), .B(_544_), .C(_558_), .Y(_487__4_) );
NOR3X1 NOR3X1_5 ( .A(_495_), .B(_532_), .C(_537_), .Y(_559_) );
AND2X2 AND2X2_35 ( .A(sumador_res_1_), .B(rom1_data_4_), .Y(_560_) );
NAND2X1 NAND2X1_81 ( .A(_560_), .B(_834_), .Y(_561_) );
INVX1 INVX1_157 ( .A(_561_), .Y(_562_) );
OAI21X1 OAI21X1_46 ( .A(_507_), .B(_530_), .C(_522_), .Y(_563_) );
NAND2X1 NAND2X1_82 ( .A(sumador_res_0_), .B(1'b0), .Y(_564_) );
INVX1 INVX1_158 ( .A(_564_), .Y(_565_) );
AND2X2 AND2X2_36 ( .A(sumador_res_2_), .B(rom1_data_3_), .Y(_566_) );
NAND2X1 NAND2X1_83 ( .A(_560_), .B(_566_), .Y(_567_) );
INVX1 INVX1_159 ( .A(rom1_data_3_), .Y(_568_) );
OAI21X1 OAI21X1_47 ( .A(_841_), .B(_568_), .C(_503_), .Y(_569_) );
NAND3X1 NAND3X1_171 ( .A(_569_), .B(_565_), .C(_567_), .Y(_570_) );
OAI21X1 OAI21X1_48 ( .A(_795_), .B(_504_), .C(_566_), .Y(_571_) );
OAI21X1 OAI21X1_49 ( .A(_841_), .B(_568_), .C(_560_), .Y(_572_) );
NAND3X1 NAND3X1_172 ( .A(_564_), .B(_571_), .C(_572_), .Y(_573_) );
AOI22X1 AOI22X1_21 ( .A(_839_), .B(_512_), .C(_516_), .D(_511_), .Y(_574_) );
NAND2X1 NAND2X1_84 ( .A(rom1_data_2_), .B(sumador_res_3_), .Y(_575_) );
INVX1 INVX1_160 ( .A(_575_), .Y(_576_) );
AND2X2 AND2X2_37 ( .A(rom1_data_0_bF_buf0_), .B(sumador_res_5_), .Y(_577_) );
NAND2X1 NAND2X1_85 ( .A(_512_), .B(_577_), .Y(_578_) );
INVX1 INVX1_161 ( .A(sumador_res_5_), .Y(_579_) );
NAND2X1 NAND2X1_86 ( .A(rom1_data_1_), .B(sumador_res_4_), .Y(_580_) );
OAI21X1 OAI21X1_50 ( .A(_777_), .B(_579_), .C(_580_), .Y(_581_) );
NAND3X1 NAND3X1_173 ( .A(_576_), .B(_581_), .C(_578_), .Y(_582_) );
NAND3X1 NAND3X1_174 ( .A(rom1_data_0_bF_buf3_), .B(sumador_res_5_), .C(_580_), .Y(_583_) );
NAND2X1 NAND2X1_87 ( .A(rom1_data_0_bF_buf2_), .B(sumador_res_5_), .Y(_584_) );
NAND3X1 NAND3X1_175 ( .A(rom1_data_1_), .B(sumador_res_4_), .C(_584_), .Y(_585_) );
NAND3X1 NAND3X1_176 ( .A(_575_), .B(_583_), .C(_585_), .Y(_586_) );
NAND3X1 NAND3X1_177 ( .A(_574_), .B(_586_), .C(_582_), .Y(_587_) );
AOI22X1 AOI22X1_22 ( .A(rom1_data_0_bF_buf1_), .B(sumador_res_4_), .C(rom1_data_1_), .D(sumador_res_3_), .Y(_588_) );
OAI22X1 OAI22X1_50 ( .A(_842_), .B(_580_), .C(_510_), .D(_588_), .Y(_589_) );
NAND3X1 NAND3X1_178 ( .A(_575_), .B(_581_), .C(_578_), .Y(_590_) );
NAND3X1 NAND3X1_179 ( .A(_576_), .B(_583_), .C(_585_), .Y(_591_) );
NAND3X1 NAND3X1_180 ( .A(_589_), .B(_591_), .C(_590_), .Y(_592_) );
AOI22X1 AOI22X1_23 ( .A(_570_), .B(_573_), .C(_587_), .D(_592_), .Y(_593_) );
NAND3X1 NAND3X1_181 ( .A(_564_), .B(_569_), .C(_567_), .Y(_594_) );
NAND3X1 NAND3X1_182 ( .A(_565_), .B(_571_), .C(_572_), .Y(_595_) );
NAND3X1 NAND3X1_183 ( .A(_589_), .B(_586_), .C(_582_), .Y(_596_) );
NAND3X1 NAND3X1_184 ( .A(_574_), .B(_591_), .C(_590_), .Y(_597_) );
AOI22X1 AOI22X1_24 ( .A(_594_), .B(_595_), .C(_596_), .D(_597_), .Y(_598_) );
OAI21X1 OAI21X1_51 ( .A(_593_), .B(_598_), .C(_563_), .Y(_599_) );
AOI21X1 AOI21X1_20 ( .A(_528_), .B(_526_), .C(_529_), .Y(_600_) );
NAND2X1 NAND2X1_88 ( .A(_570_), .B(_573_), .Y(_601_) );
AOI21X1 AOI21X1_21 ( .A(_587_), .B(_592_), .C(_601_), .Y(_602_) );
NAND2X1 NAND2X1_89 ( .A(_594_), .B(_595_), .Y(_603_) );
AOI21X1 AOI21X1_22 ( .A(_596_), .B(_597_), .C(_603_), .Y(_604_) );
OAI21X1 OAI21X1_52 ( .A(_604_), .B(_602_), .C(_600_), .Y(_605_) );
NAND3X1 NAND3X1_185 ( .A(_562_), .B(_599_), .C(_605_), .Y(_606_) );
OAI21X1 OAI21X1_53 ( .A(_593_), .B(_598_), .C(_600_), .Y(_607_) );
OAI21X1 OAI21X1_54 ( .A(_604_), .B(_602_), .C(_563_), .Y(_608_) );
NAND3X1 NAND3X1_186 ( .A(_561_), .B(_607_), .C(_608_), .Y(_609_) );
NAND3X1 NAND3X1_187 ( .A(_532_), .B(_606_), .C(_609_), .Y(_610_) );
NAND3X1 NAND3X1_188 ( .A(_561_), .B(_599_), .C(_605_), .Y(_611_) );
NAND3X1 NAND3X1_189 ( .A(_562_), .B(_607_), .C(_608_), .Y(_612_) );
NAND3X1 NAND3X1_190 ( .A(_539_), .B(_611_), .C(_612_), .Y(_613_) );
NAND3X1 NAND3X1_191 ( .A(_559_), .B(_610_), .C(_613_), .Y(_614_) );
NAND3X1 NAND3X1_192 ( .A(_539_), .B(_606_), .C(_609_), .Y(_615_) );
NAND3X1 NAND3X1_193 ( .A(_532_), .B(_611_), .C(_612_), .Y(_616_) );
NAND3X1 NAND3X1_194 ( .A(_543_), .B(_615_), .C(_616_), .Y(_617_) );
NAND2X1 NAND2X1_90 ( .A(_614_), .B(_617_), .Y(_618_) );
OAI21X1 OAI21X1_55 ( .A(_556_), .B(_554_), .C(_549_), .Y(_619_) );
NAND3X1 NAND3X1_195 ( .A(mac1_dataout_5_), .B(_614_), .C(_617_), .Y(_620_) );
INVX1 INVX1_162 ( .A(mac1_dataout_5_), .Y(_621_) );
NAND2X1 NAND2X1_91 ( .A(_621_), .B(_618_), .Y(_622_) );
NAND3X1 NAND3X1_196 ( .A(_620_), .B(_622_), .C(_619_), .Y(_623_) );
AOI21X1 AOI21X1_23 ( .A(_548_), .B(_551_), .C(_555_), .Y(_624_) );
INVX1 INVX1_163 ( .A(_620_), .Y(_625_) );
AOI21X1 AOI21X1_24 ( .A(_614_), .B(_617_), .C(mac1_dataout_5_), .Y(_626_) );
OAI21X1 OAI21X1_56 ( .A(_626_), .B(_625_), .C(_624_), .Y(_627_) );
NAND3X1 NAND3X1_197 ( .A(_745_), .B(_623_), .C(_627_), .Y(_628_) );
OAI21X1 OAI21X1_57 ( .A(_745_), .B(_618_), .C(_628_), .Y(_487__5_) );
AOI21X1 AOI21X1_25 ( .A(_615_), .B(_616_), .C(_543_), .Y(_629_) );
AOI21X1 AOI21X1_26 ( .A(_612_), .B(_611_), .C(_539_), .Y(_630_) );
NAND3X1 NAND3X1_198 ( .A(_596_), .B(_597_), .C(_603_), .Y(_631_) );
AOI21X1 AOI21X1_27 ( .A(_590_), .B(_591_), .C(_574_), .Y(_632_) );
AOI21X1 AOI21X1_28 ( .A(_582_), .B(_586_), .C(_589_), .Y(_633_) );
OAI21X1 OAI21X1_58 ( .A(_632_), .B(_633_), .C(_601_), .Y(_634_) );
AOI21X1 AOI21X1_29 ( .A(_634_), .B(_631_), .C(_563_), .Y(_635_) );
OAI21X1 OAI21X1_59 ( .A(_561_), .B(_635_), .C(_599_), .Y(_636_) );
AND2X2 AND2X2_38 ( .A(sumador_res_0_), .B(1'b0), .Y(_637_) );
NAND2X1 NAND2X1_92 ( .A(sumador_res_2_), .B(rom1_data_4_), .Y(_638_) );
OAI21X1 OAI21X1_60 ( .A(_505_), .B(_638_), .C(_570_), .Y(_639_) );
XNOR2X1 XNOR2X1_1 ( .A(_639_), .B(_637_), .Y(_640_) );
INVX1 INVX1_164 ( .A(_640_), .Y(_641_) );
OAI21X1 OAI21X1_61 ( .A(_601_), .B(_633_), .C(_596_), .Y(_642_) );
INVX1 INVX1_165 ( .A(1'b0), .Y(_643_) );
NOR2X1 NOR2X1_69 ( .A(_795_), .B(_643_), .Y(_644_) );
NAND2X1 NAND2X1_93 ( .A(sumador_res_3_), .B(rom1_data_3_), .Y(_645_) );
XOR2X1 XOR2X1_4 ( .A(_638_), .B(_645_), .Y(_646_) );
NAND2X1 NAND2X1_94 ( .A(_644_), .B(_646_), .Y(_647_) );
INVX1 INVX1_166 ( .A(_566_), .Y(_648_) );
NAND2X1 NAND2X1_95 ( .A(sumador_res_3_), .B(rom1_data_4_), .Y(_649_) );
OAI21X1 OAI21X1_62 ( .A(_846_), .B(_568_), .C(_638_), .Y(_650_) );
OAI21X1 OAI21X1_63 ( .A(_649_), .B(_648_), .C(_650_), .Y(_651_) );
OAI21X1 OAI21X1_64 ( .A(_795_), .B(_643_), .C(_651_), .Y(_652_) );
NOR2X1 NOR2X1_70 ( .A(_580_), .B(_584_), .Y(_653_) );
AOI21X1 AOI21X1_30 ( .A(_576_), .B(_581_), .C(_653_), .Y(_654_) );
NAND2X1 NAND2X1_96 ( .A(rom1_data_2_), .B(sumador_res_4_), .Y(_655_) );
INVX1 INVX1_167 ( .A(_655_), .Y(_656_) );
NAND3X1 NAND3X1_199 ( .A(rom1_data_1_), .B(sumador_res_6_), .C(_577_), .Y(_657_) );
AOI22X1 AOI22X1_25 ( .A(rom1_data_0_bF_buf0_), .B(sumador_res_6_), .C(rom1_data_1_), .D(sumador_res_5_), .Y(_658_) );
INVX1 INVX1_168 ( .A(_658_), .Y(_659_) );
NAND3X1 NAND3X1_200 ( .A(_659_), .B(_656_), .C(_657_), .Y(_660_) );
NAND2X1 NAND2X1_97 ( .A(rom1_data_1_), .B(sumador_res_6_), .Y(_661_) );
NOR2X1 NOR2X1_71 ( .A(_584_), .B(_661_), .Y(_662_) );
OAI21X1 OAI21X1_65 ( .A(_658_), .B(_662_), .C(_655_), .Y(_663_) );
NAND3X1 NAND3X1_201 ( .A(_660_), .B(_663_), .C(_654_), .Y(_664_) );
AND2X2 AND2X2_39 ( .A(_580_), .B(_584_), .Y(_665_) );
OAI21X1 OAI21X1_66 ( .A(_575_), .B(_665_), .C(_578_), .Y(_666_) );
NAND3X1 NAND3X1_202 ( .A(_655_), .B(_659_), .C(_657_), .Y(_667_) );
OAI21X1 OAI21X1_67 ( .A(_658_), .B(_662_), .C(_656_), .Y(_668_) );
NAND3X1 NAND3X1_203 ( .A(_667_), .B(_668_), .C(_666_), .Y(_669_) );
AOI22X1 AOI22X1_26 ( .A(_647_), .B(_652_), .C(_664_), .D(_669_), .Y(_670_) );
OAI21X1 OAI21X1_68 ( .A(_795_), .B(_643_), .C(_646_), .Y(_671_) );
NAND2X1 NAND2X1_98 ( .A(_644_), .B(_651_), .Y(_672_) );
NAND3X1 NAND3X1_204 ( .A(_660_), .B(_663_), .C(_666_), .Y(_673_) );
NAND3X1 NAND3X1_205 ( .A(_667_), .B(_668_), .C(_654_), .Y(_674_) );
AOI22X1 AOI22X1_27 ( .A(_671_), .B(_672_), .C(_674_), .D(_673_), .Y(_675_) );
OAI21X1 OAI21X1_69 ( .A(_670_), .B(_675_), .C(_642_), .Y(_676_) );
AOI21X1 AOI21X1_31 ( .A(_603_), .B(_597_), .C(_632_), .Y(_677_) );
AOI22X1 AOI22X1_28 ( .A(_671_), .B(_672_), .C(_664_), .D(_669_), .Y(_678_) );
AOI22X1 AOI22X1_29 ( .A(_647_), .B(_652_), .C(_674_), .D(_673_), .Y(_679_) );
OAI21X1 OAI21X1_70 ( .A(_678_), .B(_679_), .C(_677_), .Y(_680_) );
NAND3X1 NAND3X1_206 ( .A(_676_), .B(_641_), .C(_680_), .Y(_681_) );
OAI21X1 OAI21X1_71 ( .A(_670_), .B(_675_), .C(_677_), .Y(_682_) );
OAI21X1 OAI21X1_72 ( .A(_678_), .B(_679_), .C(_642_), .Y(_683_) );
NAND3X1 NAND3X1_207 ( .A(_640_), .B(_682_), .C(_683_), .Y(_684_) );
NAND3X1 NAND3X1_208 ( .A(_684_), .B(_681_), .C(_636_), .Y(_685_) );
NAND3X1 NAND3X1_209 ( .A(_596_), .B(_601_), .C(_597_), .Y(_686_) );
OAI21X1 OAI21X1_73 ( .A(_632_), .B(_633_), .C(_603_), .Y(_687_) );
AOI21X1 AOI21X1_32 ( .A(_687_), .B(_686_), .C(_600_), .Y(_688_) );
AOI21X1 AOI21X1_33 ( .A(_562_), .B(_605_), .C(_688_), .Y(_689_) );
NAND3X1 NAND3X1_210 ( .A(_640_), .B(_676_), .C(_680_), .Y(_690_) );
NAND3X1 NAND3X1_211 ( .A(_682_), .B(_641_), .C(_683_), .Y(_691_) );
NAND3X1 NAND3X1_212 ( .A(_690_), .B(_691_), .C(_689_), .Y(_692_) );
NAND3X1 NAND3X1_213 ( .A(_630_), .B(_692_), .C(_685_), .Y(_693_) );
NAND3X1 NAND3X1_214 ( .A(_684_), .B(_681_), .C(_689_), .Y(_694_) );
NAND3X1 NAND3X1_215 ( .A(_690_), .B(_691_), .C(_636_), .Y(_695_) );
NAND3X1 NAND3X1_216 ( .A(_610_), .B(_694_), .C(_695_), .Y(_696_) );
NAND3X1 NAND3X1_217 ( .A(_629_), .B(_693_), .C(_696_), .Y(_697_) );
NAND3X1 NAND3X1_218 ( .A(_610_), .B(_692_), .C(_685_), .Y(_698_) );
NAND3X1 NAND3X1_219 ( .A(_630_), .B(_694_), .C(_695_), .Y(_699_) );
NAND3X1 NAND3X1_220 ( .A(_614_), .B(_698_), .C(_699_), .Y(_700_) );
NAND2X1 NAND2X1_99 ( .A(_697_), .B(_700_), .Y(_701_) );
OAI21X1 OAI21X1_74 ( .A(_626_), .B(_624_), .C(_620_), .Y(_702_) );
NAND3X1 NAND3X1_221 ( .A(mac1_dataout_6_), .B(_697_), .C(_700_), .Y(_703_) );
INVX1 INVX1_169 ( .A(mac1_dataout_6_), .Y(_704_) );
NAND3X1 NAND3X1_222 ( .A(_614_), .B(_693_), .C(_696_), .Y(_705_) );
NAND3X1 NAND3X1_223 ( .A(_629_), .B(_698_), .C(_699_), .Y(_706_) );
NAND3X1 NAND3X1_224 ( .A(_704_), .B(_705_), .C(_706_), .Y(_707_) );
AOI21X1 AOI21X1_34 ( .A(_703_), .B(_707_), .C(_702_), .Y(_708_) );
AOI21X1 AOI21X1_35 ( .A(_619_), .B(_622_), .C(_625_), .Y(_709_) );
NAND2X1 NAND2X1_100 ( .A(_703_), .B(_707_), .Y(_710_) );
OAI21X1 OAI21X1_75 ( .A(_709_), .B(_710_), .C(_745_), .Y(_711_) );
OAI22X1 OAI22X1_51 ( .A(_745_), .B(_701_), .C(_708_), .D(_711_), .Y(_487__6_) );
NAND2X1 NAND2X1_101 ( .A(_693_), .B(_697_), .Y(_712_) );
INVX1 INVX1_170 ( .A(_712_), .Y(_713_) );
INVX1 INVX1_171 ( .A(_685_), .Y(_714_) );
NAND2X1 NAND2X1_102 ( .A(_637_), .B(_639_), .Y(_715_) );
INVX1 INVX1_172 ( .A(_715_), .Y(_716_) );
NAND2X1 NAND2X1_103 ( .A(_676_), .B(_681_), .Y(_717_) );
OAI21X1 OAI21X1_76 ( .A(_648_), .B(_649_), .C(_647_), .Y(_718_) );
NAND2X1 NAND2X1_104 ( .A(sumador_res_0_), .B(1'b0), .Y(_719_) );
NAND2X1 NAND2X1_105 ( .A(sumador_res_1_), .B(1'b0), .Y(_720_) );
XOR2X1 XOR2X1_5 ( .A(_719_), .B(_720_), .Y(_721_) );
XOR2X1 XOR2X1_6 ( .A(_718_), .B(_721_), .Y(_722_) );
INVX1 INVX1_173 ( .A(_722_), .Y(_723_) );
INVX1 INVX1_174 ( .A(_673_), .Y(_724_) );
OR2X2 OR2X2_3 ( .A(_678_), .B(_724_), .Y(_725_) );
INVX1 INVX1_175 ( .A(rom1_data_2_), .Y(_726_) );
NOR2X1 NOR2X1_72 ( .A(_726_), .B(_579_), .Y(_727_) );
NAND2X1 NAND2X1_106 ( .A(rom1_data_0_bF_buf3_), .B(sumador_res_7_), .Y(_728_) );
XNOR2X1 XNOR2X1_2 ( .A(_661_), .B(_728_), .Y(_729_) );
INVX1 INVX1_176 ( .A(_729_), .Y(_730_) );
NAND2X1 NAND2X1_107 ( .A(_727_), .B(_730_), .Y(_731_) );
OAI21X1 OAI21X1_77 ( .A(_726_), .B(_579_), .C(_729_), .Y(_732_) );
OAI21X1 OAI21X1_78 ( .A(_655_), .B(_658_), .C(_657_), .Y(_733_) );
INVX1 INVX1_177 ( .A(_733_), .Y(_735_) );
NAND3X1 NAND3X1_225 ( .A(_732_), .B(_735_), .C(_731_), .Y(_736_) );
NAND2X1 NAND2X1_108 ( .A(_727_), .B(_729_), .Y(_737_) );
OAI21X1 OAI21X1_79 ( .A(_726_), .B(_579_), .C(_730_), .Y(_738_) );
NAND3X1 NAND3X1_226 ( .A(_733_), .B(_737_), .C(_738_), .Y(_739_) );
NAND2X1 NAND2X1_109 ( .A(rom1_data_3_), .B(sumador_res_4_), .Y(_740_) );
XNOR2X1 XNOR2X1_3 ( .A(_649_), .B(_740_), .Y(_741_) );
NAND2X1 NAND2X1_110 ( .A(sumador_res_2_), .B(1'b0), .Y(_742_) );
XOR2X1 XOR2X1_7 ( .A(_741_), .B(_742_), .Y(_743_) );
INVX1 INVX1_178 ( .A(_743_), .Y(_744_) );
NAND3X1 NAND3X1_227 ( .A(_736_), .B(_739_), .C(_744_), .Y(_746_) );
NAND3X1 NAND3X1_228 ( .A(_732_), .B(_733_), .C(_731_), .Y(_747_) );
NAND3X1 NAND3X1_229 ( .A(_735_), .B(_737_), .C(_738_), .Y(_748_) );
NAND3X1 NAND3X1_230 ( .A(_743_), .B(_747_), .C(_748_), .Y(_749_) );
NAND3X1 NAND3X1_231 ( .A(_749_), .B(_746_), .C(_725_), .Y(_750_) );
NOR2X1 NOR2X1_73 ( .A(_724_), .B(_678_), .Y(_751_) );
NAND3X1 NAND3X1_232 ( .A(_747_), .B(_748_), .C(_744_), .Y(_752_) );
NAND3X1 NAND3X1_233 ( .A(_743_), .B(_736_), .C(_739_), .Y(_753_) );
NAND3X1 NAND3X1_234 ( .A(_751_), .B(_753_), .C(_752_), .Y(_754_) );
AOI21X1 AOI21X1_36 ( .A(_750_), .B(_754_), .C(_723_), .Y(_755_) );
NAND3X1 NAND3X1_235 ( .A(_751_), .B(_749_), .C(_746_), .Y(_757_) );
NAND3X1 NAND3X1_236 ( .A(_753_), .B(_752_), .C(_725_), .Y(_758_) );
AOI21X1 AOI21X1_37 ( .A(_758_), .B(_757_), .C(_722_), .Y(_759_) );
OAI21X1 OAI21X1_80 ( .A(_755_), .B(_759_), .C(_717_), .Y(_760_) );
INVX1 INVX1_179 ( .A(_717_), .Y(_761_) );
NAND3X1 NAND3X1_237 ( .A(_722_), .B(_757_), .C(_758_), .Y(_762_) );
NAND3X1 NAND3X1_238 ( .A(_723_), .B(_754_), .C(_750_), .Y(_763_) );
NAND3X1 NAND3X1_239 ( .A(_762_), .B(_763_), .C(_761_), .Y(_764_) );
AOI21X1 AOI21X1_38 ( .A(_764_), .B(_760_), .C(_716_), .Y(_765_) );
NAND3X1 NAND3X1_240 ( .A(_717_), .B(_762_), .C(_763_), .Y(_766_) );
OAI21X1 OAI21X1_81 ( .A(_755_), .B(_759_), .C(_761_), .Y(_767_) );
AOI21X1 AOI21X1_39 ( .A(_767_), .B(_766_), .C(_715_), .Y(_768_) );
OAI21X1 OAI21X1_82 ( .A(_768_), .B(_765_), .C(_714_), .Y(_769_) );
NAND3X1 NAND3X1_241 ( .A(_715_), .B(_766_), .C(_767_), .Y(_770_) );
NAND3X1 NAND3X1_242 ( .A(_716_), .B(_760_), .C(_764_), .Y(_771_) );
NAND3X1 NAND3X1_243 ( .A(_685_), .B(_770_), .C(_771_), .Y(_772_) );
NAND3X1 NAND3X1_244 ( .A(_713_), .B(_772_), .C(_769_), .Y(_773_) );
NAND2X1 NAND2X1_111 ( .A(_760_), .B(_764_), .Y(_774_) );
XOR2X1 XOR2X1_8 ( .A(_685_), .B(_716_), .Y(_775_) );
OR2X2 OR2X2_4 ( .A(_774_), .B(_775_), .Y(_776_) );
NAND2X1 NAND2X1_112 ( .A(_775_), .B(_774_), .Y(_778_) );
NAND3X1 NAND3X1_245 ( .A(_712_), .B(_778_), .C(_776_), .Y(_779_) );
NAND2X1 NAND2X1_113 ( .A(_779_), .B(_773_), .Y(_780_) );
INVX1 INVX1_180 ( .A(mac1_dataout_7_), .Y(_781_) );
AOI21X1 AOI21X1_40 ( .A(_705_), .B(_706_), .C(_704_), .Y(_782_) );
AOI21X1 AOI21X1_41 ( .A(_702_), .B(_707_), .C(_782_), .Y(_783_) );
NAND2X1 NAND2X1_114 ( .A(_781_), .B(_783_), .Y(_784_) );
AOI21X1 AOI21X1_42 ( .A(_697_), .B(_700_), .C(mac1_dataout_6_), .Y(_785_) );
OAI21X1 OAI21X1_83 ( .A(_785_), .B(_709_), .C(_703_), .Y(_786_) );
AOI21X1 AOI21X1_43 ( .A(_786_), .B(mac1_dataout_7_), .C(mac1_reset_bF_buf0), .Y(_787_) );
NAND3X1 NAND3X1_246 ( .A(_780_), .B(_784_), .C(_787_), .Y(_789_) );
AOI21X1 AOI21X1_44 ( .A(_776_), .B(_778_), .C(_713_), .Y(_790_) );
AOI21X1 AOI21X1_45 ( .A(_769_), .B(_772_), .C(_712_), .Y(_791_) );
AND2X2 AND2X2_40 ( .A(_783_), .B(_781_), .Y(_792_) );
OAI21X1 OAI21X1_84 ( .A(_781_), .B(_783_), .C(_745_), .Y(_793_) );
OAI22X1 OAI22X1_52 ( .A(_790_), .B(_791_), .C(_793_), .D(_792_), .Y(_794_) );
NAND2X1 NAND2X1_115 ( .A(_794_), .B(_789_), .Y(_487__7_) );
DFFPOSX1 DFFPOSX1_14 ( .CLK(clk_bF_buf2), .D(_487__0_), .Q(mac1_dataout_0_) );
DFFPOSX1 DFFPOSX1_15 ( .CLK(clk_bF_buf2), .D(_487__1_), .Q(mac1_dataout_1_) );
DFFPOSX1 DFFPOSX1_16 ( .CLK(clk_bF_buf5), .D(_487__2_), .Q(mac1_dataout_2_) );
DFFPOSX1 DFFPOSX1_17 ( .CLK(clk_bF_buf1), .D(_487__3_), .Q(mac1_dataout_3_) );
DFFPOSX1 DFFPOSX1_18 ( .CLK(clk_bF_buf0), .D(_487__4_), .Q(mac1_dataout_4_) );
DFFPOSX1 DFFPOSX1_19 ( .CLK(clk_bF_buf5), .D(_487__5_), .Q(mac1_dataout_5_) );
DFFPOSX1 DFFPOSX1_20 ( .CLK(clk_bF_buf2), .D(_487__6_), .Q(mac1_dataout_6_) );
DFFPOSX1 DFFPOSX1_21 ( .CLK(clk_bF_buf3), .D(_487__7_), .Q(mac1_dataout_7_) );
INVX1 INVX1_181 ( .A(reg1_dataout_0_), .Y(_855_) );
NAND2X1 NAND2X1_116 ( .A(din[0]), .B(1'b1), .Y(_856_) );
OAI21X1 OAI21X1_85 ( .A(1'b1), .B(_855_), .C(_856_), .Y(_853__0_) );
INVX1 INVX1_182 ( .A(reg1_dataout_1_), .Y(_857_) );
NAND2X1 NAND2X1_117 ( .A(1'b1), .B(din[1]), .Y(_858_) );
OAI21X1 OAI21X1_86 ( .A(1'b1), .B(_857_), .C(_858_), .Y(_853__1_) );
INVX1 INVX1_183 ( .A(reg1_dataout_2_), .Y(_859_) );
NAND2X1 NAND2X1_118 ( .A(1'b1), .B(din[2]), .Y(_860_) );
OAI21X1 OAI21X1_87 ( .A(1'b1), .B(_859_), .C(_860_), .Y(_853__2_) );
INVX1 INVX1_184 ( .A(reg1_dataout_3_), .Y(_861_) );
NAND2X1 NAND2X1_119 ( .A(1'b1), .B(din[3]), .Y(_862_) );
OAI21X1 OAI21X1_88 ( .A(1'b1), .B(_861_), .C(_862_), .Y(_853__3_) );
INVX1 INVX1_185 ( .A(reg1_dataout_4_), .Y(_863_) );
NAND2X1 NAND2X1_120 ( .A(1'b1), .B(din[4]), .Y(_864_) );
OAI21X1 OAI21X1_89 ( .A(1'b1), .B(_863_), .C(_864_), .Y(_853__4_) );
INVX1 INVX1_186 ( .A(reg1_dataout_5_), .Y(_865_) );
NAND2X1 NAND2X1_121 ( .A(1'b1), .B(din[5]), .Y(_866_) );
OAI21X1 OAI21X1_90 ( .A(1'b1), .B(_865_), .C(_866_), .Y(_853__5_) );
INVX1 INVX1_187 ( .A(reg1_dataout_6_), .Y(_867_) );
NAND2X1 NAND2X1_122 ( .A(1'b1), .B(din[6]), .Y(_868_) );
OAI21X1 OAI21X1_91 ( .A(1'b1), .B(_867_), .C(_868_), .Y(_853__6_) );
INVX1 INVX1_188 ( .A(reg1_dataout_7_), .Y(_869_) );
NAND2X1 NAND2X1_123 ( .A(1'b1), .B(din[7]), .Y(_870_) );
OAI21X1 OAI21X1_92 ( .A(1'b1), .B(_869_), .C(_870_), .Y(_853__7_) );
INVX1 INVX1_189 ( .A(rst_bF_buf3), .Y(_854_) );
DFFSR DFFSR_257 ( .CLK(clk2_clkout_bF_buf23), .D(_853__0_), .Q(reg1_dataout_0_), .R(_854_), .S(1'b1) );
DFFSR DFFSR_258 ( .CLK(clk2_clkout_bF_buf38), .D(_853__1_), .Q(reg1_dataout_1_), .R(_854_), .S(1'b1) );
DFFSR DFFSR_259 ( .CLK(clk2_clkout_bF_buf41), .D(_853__2_), .Q(reg1_dataout_2_), .R(_854_), .S(1'b1) );
DFFSR DFFSR_260 ( .CLK(clk2_clkout_bF_buf38), .D(_853__3_), .Q(reg1_dataout_3_), .R(_854_), .S(1'b1) );
DFFSR DFFSR_261 ( .CLK(clk2_clkout_bF_buf12), .D(_853__4_), .Q(reg1_dataout_4_), .R(_854_), .S(1'b1) );
DFFSR DFFSR_262 ( .CLK(clk2_clkout_bF_buf14), .D(_853__5_), .Q(reg1_dataout_5_), .R(_854_), .S(1'b1) );
DFFSR DFFSR_263 ( .CLK(clk2_clkout_bF_buf34), .D(_853__6_), .Q(reg1_dataout_6_), .R(_854_), .S(1'b1) );
DFFSR DFFSR_264 ( .CLK(clk2_clkout_bF_buf38), .D(_853__7_), .Q(reg1_dataout_7_), .R(_854_), .S(1'b1) );
INVX1 INVX1_190 ( .A(reg2_dataout_0_), .Y(_873_) );
NAND2X1 NAND2X1_124 ( .A(mac1_dataout_0_), .B(mac1_reset_bF_buf1), .Y(_874_) );
OAI21X1 OAI21X1_93 ( .A(mac1_reset_bF_buf1), .B(_873_), .C(_874_), .Y(_871__0_) );
INVX1 INVX1_191 ( .A(reg2_dataout_1_), .Y(_875_) );
NAND2X1 NAND2X1_125 ( .A(mac1_reset_bF_buf1), .B(mac1_dataout_1_), .Y(_876_) );
OAI21X1 OAI21X1_94 ( .A(mac1_reset_bF_buf1), .B(_875_), .C(_876_), .Y(_871__1_) );
INVX1 INVX1_192 ( .A(reg2_dataout_2_), .Y(_877_) );
NAND2X1 NAND2X1_126 ( .A(mac1_reset_bF_buf2), .B(mac1_dataout_2_), .Y(_878_) );
OAI21X1 OAI21X1_95 ( .A(mac1_reset_bF_buf2), .B(_877_), .C(_878_), .Y(_871__2_) );
INVX1 INVX1_193 ( .A(reg2_dataout_3_), .Y(_879_) );
NAND2X1 NAND2X1_127 ( .A(mac1_reset_bF_buf0), .B(mac1_dataout_3_), .Y(_880_) );
OAI21X1 OAI21X1_96 ( .A(mac1_reset_bF_buf0), .B(_879_), .C(_880_), .Y(_871__3_) );
INVX1 INVX1_194 ( .A(reg2_dataout_4_), .Y(_881_) );
NAND2X1 NAND2X1_128 ( .A(mac1_reset_bF_buf2), .B(mac1_dataout_4_), .Y(_882_) );
OAI21X1 OAI21X1_97 ( .A(mac1_reset_bF_buf2), .B(_881_), .C(_882_), .Y(_871__4_) );
INVX1 INVX1_195 ( .A(reg2_dataout_5_), .Y(_883_) );
NAND2X1 NAND2X1_129 ( .A(mac1_reset_bF_buf3), .B(mac1_dataout_5_), .Y(_884_) );
OAI21X1 OAI21X1_98 ( .A(mac1_reset_bF_buf3), .B(_883_), .C(_884_), .Y(_871__5_) );
INVX1 INVX1_196 ( .A(reg2_dataout_6_), .Y(_885_) );
NAND2X1 NAND2X1_130 ( .A(mac1_reset_bF_buf3), .B(mac1_dataout_6_), .Y(_886_) );
OAI21X1 OAI21X1_99 ( .A(mac1_reset_bF_buf3), .B(_885_), .C(_886_), .Y(_871__6_) );
INVX1 INVX1_197 ( .A(reg2_dataout_7_), .Y(_887_) );
NAND2X1 NAND2X1_131 ( .A(mac1_reset_bF_buf0), .B(mac1_dataout_7_), .Y(_888_) );
OAI21X1 OAI21X1_100 ( .A(mac1_reset_bF_buf0), .B(_887_), .C(_888_), .Y(_871__7_) );
INVX1 INVX1_198 ( .A(rst_bF_buf2), .Y(_872_) );
DFFSR DFFSR_265 ( .CLK(clk_bF_buf2), .D(_871__0_), .Q(reg2_dataout_0_), .R(_872_), .S(1'b1) );
DFFSR DFFSR_266 ( .CLK(clk_bF_buf2), .D(_871__1_), .Q(reg2_dataout_1_), .R(_872_), .S(1'b1) );
DFFSR DFFSR_267 ( .CLK(clk_bF_buf5), .D(_871__2_), .Q(reg2_dataout_2_), .R(_872_), .S(1'b1) );
DFFSR DFFSR_268 ( .CLK(clk_bF_buf1), .D(_871__3_), .Q(reg2_dataout_3_), .R(_872_), .S(1'b1) );
DFFSR DFFSR_269 ( .CLK(clk_bF_buf2), .D(_871__4_), .Q(reg2_dataout_4_), .R(_872_), .S(1'b1) );
DFFSR DFFSR_270 ( .CLK(clk_bF_buf5), .D(_871__5_), .Q(reg2_dataout_5_), .R(_872_), .S(1'b1) );
DFFSR DFFSR_271 ( .CLK(clk_bF_buf1), .D(_871__6_), .Q(reg2_dataout_6_), .R(_872_), .S(1'b1) );
DFFSR DFFSR_272 ( .CLK(clk_bF_buf4), .D(_871__7_), .Q(reg2_dataout_7_), .R(_872_), .S(1'b1) );
INVX1 INVX1_199 ( .A(reg3_dataout_0_), .Y(_891_) );
NAND2X1 NAND2X1_132 ( .A(reg2_dataout_0_), .B(1'b1), .Y(_892_) );
OAI21X1 OAI21X1_101 ( .A(1'b1), .B(_891_), .C(_892_), .Y(_889__0_) );
INVX1 INVX1_200 ( .A(reg3_dataout_1_), .Y(_893_) );
NAND2X1 NAND2X1_133 ( .A(1'b1), .B(reg2_dataout_1_), .Y(_894_) );
OAI21X1 OAI21X1_102 ( .A(1'b1), .B(_893_), .C(_894_), .Y(_889__1_) );
INVX1 INVX1_201 ( .A(reg3_dataout_2_), .Y(_895_) );
NAND2X1 NAND2X1_134 ( .A(1'b1), .B(reg2_dataout_2_), .Y(_896_) );
OAI21X1 OAI21X1_103 ( .A(1'b1), .B(_895_), .C(_896_), .Y(_889__2_) );
INVX1 INVX1_202 ( .A(reg3_dataout_3_), .Y(_897_) );
NAND2X1 NAND2X1_135 ( .A(1'b1), .B(reg2_dataout_3_), .Y(_898_) );
OAI21X1 OAI21X1_104 ( .A(1'b1), .B(_897_), .C(_898_), .Y(_889__3_) );
INVX1 INVX1_203 ( .A(reg3_dataout_4_), .Y(_899_) );
NAND2X1 NAND2X1_136 ( .A(1'b1), .B(reg2_dataout_4_), .Y(_900_) );
OAI21X1 OAI21X1_105 ( .A(1'b1), .B(_899_), .C(_900_), .Y(_889__4_) );
INVX1 INVX1_204 ( .A(reg3_dataout_5_), .Y(_901_) );
NAND2X1 NAND2X1_137 ( .A(1'b1), .B(reg2_dataout_5_), .Y(_902_) );
OAI21X1 OAI21X1_106 ( .A(1'b1), .B(_901_), .C(_902_), .Y(_889__5_) );
INVX1 INVX1_205 ( .A(reg3_dataout_6_), .Y(_903_) );
NAND2X1 NAND2X1_138 ( .A(1'b1), .B(reg2_dataout_6_), .Y(_904_) );
OAI21X1 OAI21X1_107 ( .A(1'b1), .B(_903_), .C(_904_), .Y(_889__6_) );
INVX1 INVX1_206 ( .A(reg3_dataout_7_), .Y(_905_) );
NAND2X1 NAND2X1_139 ( .A(1'b1), .B(reg2_dataout_7_), .Y(_906_) );
OAI21X1 OAI21X1_108 ( .A(1'b1), .B(_905_), .C(_906_), .Y(_889__7_) );
INVX1 INVX1_207 ( .A(rst_bF_buf5), .Y(_890_) );
DFFSR DFFSR_273 ( .CLK(clk2_clkout_bF_buf27), .D(_889__0_), .Q(reg3_dataout_0_), .R(_890_), .S(1'b1) );
DFFSR DFFSR_274 ( .CLK(clk2_clkout_bF_buf27), .D(_889__1_), .Q(reg3_dataout_1_), .R(_890_), .S(1'b1) );
DFFSR DFFSR_275 ( .CLK(clk2_clkout_bF_buf14), .D(_889__2_), .Q(reg3_dataout_2_), .R(_890_), .S(1'b1) );
DFFSR DFFSR_276 ( .CLK(clk2_clkout_bF_buf27), .D(_889__3_), .Q(reg3_dataout_3_), .R(_890_), .S(1'b1) );
DFFSR DFFSR_277 ( .CLK(clk2_clkout_bF_buf27), .D(_889__4_), .Q(reg3_dataout_4_), .R(_890_), .S(1'b1) );
DFFSR DFFSR_278 ( .CLK(clk2_clkout_bF_buf27), .D(_889__5_), .Q(reg3_dataout_5_), .R(_890_), .S(1'b1) );
DFFSR DFFSR_279 ( .CLK(clk2_clkout_bF_buf14), .D(_889__6_), .Q(reg3_dataout_6_), .R(_890_), .S(1'b1) );
DFFSR DFFSR_280 ( .CLK(clk2_clkout_bF_buf9), .D(_889__7_), .Q(reg3_dataout_7_), .R(_890_), .S(1'b1) );
INVX1 INVX1_208 ( .A(1'b1), .Y(_923_) );
NAND2X1 NAND2X1_140 ( .A(ret2_rf_13_), .B(_923_), .Y(_924_) );
NAND2X1 NAND2X1_141 ( .A(ret2_rf_12_), .B(1'b1), .Y(_925_) );
AOI21X1 AOI21X1_46 ( .A(_924_), .B(_925_), .C(rst_bF_buf1), .Y(_912_) );
NAND2X1 NAND2X1_142 ( .A(ret2_rf_14_), .B(_923_), .Y(_926_) );
NAND2X1 NAND2X1_143 ( .A(ret2_rf_13_), .B(1'b1), .Y(_927_) );
AOI21X1 AOI21X1_47 ( .A(_926_), .B(_927_), .C(rst_bF_buf4), .Y(_913_) );
NAND2X1 NAND2X1_144 ( .A(ret2_rf_12_), .B(_923_), .Y(_928_) );
NAND2X1 NAND2X1_145 ( .A(1'b1), .B(ret2_rf_11_), .Y(_929_) );
AOI21X1 AOI21X1_48 ( .A(_928_), .B(_929_), .C(rst_bF_buf1), .Y(_911_) );
NAND2X1 NAND2X1_146 ( .A(ret2_rf_11_), .B(_923_), .Y(_930_) );
NAND2X1 NAND2X1_147 ( .A(1'b1), .B(ret2_rf_10_), .Y(_931_) );
AOI21X1 AOI21X1_49 ( .A(_930_), .B(_931_), .C(rst_bF_buf4), .Y(_910_) );
NAND2X1 NAND2X1_148 ( .A(ret2_rf_10_), .B(_923_), .Y(_932_) );
NAND2X1 NAND2X1_149 ( .A(1'b1), .B(ret2_rf_9_), .Y(_933_) );
AOI21X1 AOI21X1_50 ( .A(_932_), .B(_933_), .C(rst_bF_buf4), .Y(_909_) );
NAND2X1 NAND2X1_150 ( .A(ret2_rf_9_), .B(_923_), .Y(_934_) );
NAND2X1 NAND2X1_151 ( .A(1'b1), .B(ret2_rf_8_), .Y(_935_) );
AOI21X1 AOI21X1_51 ( .A(_934_), .B(_935_), .C(rst_bF_buf5), .Y(_922_) );
NAND2X1 NAND2X1_152 ( .A(ret2_rf_8_), .B(_923_), .Y(_936_) );
NAND2X1 NAND2X1_153 ( .A(1'b1), .B(ret2_rf_7_), .Y(_937_) );
AOI21X1 AOI21X1_52 ( .A(_936_), .B(_937_), .C(rst_bF_buf3), .Y(_921_) );
NAND2X1 NAND2X1_154 ( .A(ret2_rf_7_), .B(_923_), .Y(_938_) );
NAND2X1 NAND2X1_155 ( .A(1'b1), .B(ret2_rf_6_), .Y(_939_) );
AOI21X1 AOI21X1_53 ( .A(_938_), .B(_939_), .C(rst_bF_buf0), .Y(_920_) );
NAND2X1 NAND2X1_156 ( .A(ret2_rf_6_), .B(_923_), .Y(_940_) );
NAND2X1 NAND2X1_157 ( .A(1'b1), .B(ret2_rf_5_), .Y(_941_) );
AOI21X1 AOI21X1_54 ( .A(_940_), .B(_941_), .C(rst_bF_buf5), .Y(_919_) );
NAND2X1 NAND2X1_158 ( .A(ret2_rf_5_), .B(_923_), .Y(_942_) );
NAND2X1 NAND2X1_159 ( .A(1'b1), .B(ret2_rf_4_), .Y(_943_) );
AOI21X1 AOI21X1_55 ( .A(_942_), .B(_943_), .C(rst_bF_buf3), .Y(_918_) );
NAND2X1 NAND2X1_160 ( .A(ret2_rf_4_), .B(_923_), .Y(_944_) );
NAND2X1 NAND2X1_161 ( .A(1'b1), .B(ret2_rf_3_), .Y(_945_) );
AOI21X1 AOI21X1_56 ( .A(_944_), .B(_945_), .C(rst_bF_buf3), .Y(_917_) );
NAND2X1 NAND2X1_162 ( .A(ret2_rf_3_), .B(_923_), .Y(_946_) );
NAND2X1 NAND2X1_163 ( .A(1'b1), .B(ret2_rf_2_), .Y(_947_) );
AOI21X1 AOI21X1_57 ( .A(_946_), .B(_947_), .C(rst_bF_buf4), .Y(_916_) );
NAND2X1 NAND2X1_164 ( .A(ret2_rf_2_), .B(_923_), .Y(_948_) );
NAND2X1 NAND2X1_165 ( .A(1'b1), .B(ret2_rf_1_), .Y(_949_) );
AOI21X1 AOI21X1_58 ( .A(_948_), .B(_949_), .C(rst_bF_buf4), .Y(_915_) );
NAND2X1 NAND2X1_166 ( .A(ret2_rf_1_), .B(_923_), .Y(_950_) );
NAND2X1 NAND2X1_167 ( .A(1'b1), .B(ret2_rf_0_), .Y(_951_) );
AOI21X1 AOI21X1_59 ( .A(_950_), .B(_951_), .C(rst_bF_buf5), .Y(_914_) );
NAND2X1 NAND2X1_168 ( .A(ret2_rf_0_), .B(_923_), .Y(_952_) );
NAND2X1 NAND2X1_169 ( .A(1'b1), .B(comp_dataout), .Y(_953_) );
AOI21X1 AOI21X1_60 ( .A(_952_), .B(_953_), .C(rst_bF_buf0), .Y(_908_) );
NAND2X1 NAND2X1_170 ( .A(1'b1), .B(ret2_rf_14_), .Y(_954_) );
NOR2X1 NOR2X1_74 ( .A(rst_bF_buf1), .B(_954_), .Y(_907_) );
DFFPOSX1 DFFPOSX1_22 ( .CLK(clk_bF_buf0), .D(_907_), .Q(mac1_reset) );
DFFPOSX1 DFFPOSX1_23 ( .CLK(clk_bF_buf4), .D(_917_), .Q(ret2_rf_4_) );
DFFPOSX1 DFFPOSX1_24 ( .CLK(clk_bF_buf1), .D(_914_), .Q(ret2_rf_1_) );
DFFPOSX1 DFFPOSX1_25 ( .CLK(clk_bF_buf3), .D(_908_), .Q(ret2_rf_0_) );
DFFPOSX1 DFFPOSX1_26 ( .CLK(clk_bF_buf4), .D(_919_), .Q(ret2_rf_6_) );
DFFPOSX1 DFFPOSX1_27 ( .CLK(clk_bF_buf0), .D(_922_), .Q(ret2_rf_9_) );
DFFPOSX1 DFFPOSX1_28 ( .CLK(clk_bF_buf6), .D(_909_), .Q(ret2_rf_10_) );
DFFPOSX1 DFFPOSX1_29 ( .CLK(clk_bF_buf5), .D(_916_), .Q(ret2_rf_3_) );
DFFPOSX1 DFFPOSX1_30 ( .CLK(clk_bF_buf3), .D(_920_), .Q(ret2_rf_7_) );
DFFPOSX1 DFFPOSX1_31 ( .CLK(clk_bF_buf4), .D(_921_), .Q(ret2_rf_8_) );
DFFPOSX1 DFFPOSX1_32 ( .CLK(clk_bF_buf5), .D(_915_), .Q(ret2_rf_2_) );
DFFPOSX1 DFFPOSX1_33 ( .CLK(clk_bF_buf4), .D(_918_), .Q(ret2_rf_5_) );
DFFPOSX1 DFFPOSX1_34 ( .CLK(clk_bF_buf6), .D(_910_), .Q(ret2_rf_11_) );
DFFPOSX1 DFFPOSX1_35 ( .CLK(clk_bF_buf0), .D(_911_), .Q(ret2_rf_12_) );
DFFPOSX1 DFFPOSX1_36 ( .CLK(clk_bF_buf6), .D(_912_), .Q(ret2_rf_13_) );
DFFPOSX1 DFFPOSX1_37 ( .CLK(clk_bF_buf6), .D(_913_), .Q(ret2_rf_14_) );
NOR2X1 NOR2X1_75 ( .A(counterup_counter_0_bF_buf2_), .B(rst_bF_buf5), .Y(_955__0_) );
INVX1 INVX1_209 ( .A(rst_bF_buf3), .Y(_956_) );
OAI21X1 OAI21X1_109 ( .A(counterup_counter_0_bF_buf1_), .B(counterup_counter_1_), .C(_956_), .Y(_957_) );
AOI21X1 AOI21X1_61 ( .A(counterup_counter_0_bF_buf0_), .B(counterup_counter_1_), .C(_957_), .Y(_955__1_) );
AOI21X1 AOI21X1_62 ( .A(counterup_counter_0_bF_buf3_), .B(counterup_counter_1_), .C(counterup_counter_2_), .Y(_958_) );
NAND3X1 NAND3X1_247 ( .A(counterup_counter_0_bF_buf2_), .B(counterup_counter_1_), .C(counterup_counter_2_), .Y(_959_) );
NAND2X1 NAND2X1_171 ( .A(_956_), .B(_959_), .Y(_960_) );
NOR2X1 NOR2X1_76 ( .A(_958_), .B(_960_), .Y(_955__2_) );
INVX1 INVX1_210 ( .A(counterup_counter_3_), .Y(_961_) );
OAI21X1 OAI21X1_110 ( .A(_961_), .B(_959_), .C(_956_), .Y(_962_) );
AOI21X1 AOI21X1_63 ( .A(_961_), .B(_959_), .C(_962_), .Y(_955__3_) );
NOR3X1 NOR3X1_6 ( .A(rst_bF_buf3), .B(_961_), .C(_959_), .Y(_955__4_) );
DFFPOSX1 DFFPOSX1_38 ( .CLK(clk_bF_buf1), .D(_955__0_), .Q(rom1_data_0_) );
DFFPOSX1 DFFPOSX1_39 ( .CLK(clk_bF_buf5), .D(_955__1_), .Q(rom1_data_1_) );
DFFPOSX1 DFFPOSX1_40 ( .CLK(clk_bF_buf1), .D(_955__2_), .Q(rom1_data_2_) );
DFFPOSX1 DFFPOSX1_41 ( .CLK(clk_bF_buf3), .D(_955__3_), .Q(rom1_data_3_) );
DFFPOSX1 DFFPOSX1_42 ( .CLK(clk_bF_buf2), .D(_955__4_), .Q(rom1_data_4_) );
NAND2X1 NAND2X1_172 ( .A(asr1_dataout_0_), .B(asr2_dataout_0_), .Y(_964_) );
INVX1 INVX1_211 ( .A(_964_), .Y(_965_) );
INVX1 INVX1_212 ( .A(rst_bF_buf0), .Y(_966_) );
OAI21X1 OAI21X1_111 ( .A(asr1_dataout_0_), .B(asr2_dataout_0_), .C(_966_), .Y(_967_) );
NOR2X1 NOR2X1_77 ( .A(_965_), .B(_967_), .Y(_963__0_) );
XOR2X1 XOR2X1_9 ( .A(asr1_dataout_1_), .B(asr2_dataout_1_), .Y(_968_) );
AND2X2 AND2X2_41 ( .A(_968_), .B(_965_), .Y(_969_) );
OAI21X1 OAI21X1_112 ( .A(_965_), .B(_968_), .C(_966_), .Y(_970_) );
OR2X2 OR2X2_5 ( .A(_969_), .B(_970_), .Y(_971_) );
INVX1 INVX1_213 ( .A(_971_), .Y(_963__1_) );
NOR2X1 NOR2X1_78 ( .A(asr1_dataout_1_), .B(asr2_dataout_1_), .Y(_972_) );
NAND2X1 NAND2X1_173 ( .A(asr1_dataout_1_), .B(asr2_dataout_1_), .Y(_973_) );
OAI21X1 OAI21X1_113 ( .A(_964_), .B(_972_), .C(_973_), .Y(_974_) );
XOR2X1 XOR2X1_10 ( .A(asr1_dataout_2_), .B(asr2_dataout_2_), .Y(_975_) );
OAI21X1 OAI21X1_114 ( .A(_975_), .B(_974_), .C(_966_), .Y(_976_) );
AOI21X1 AOI21X1_64 ( .A(_974_), .B(_975_), .C(_976_), .Y(_963__2_) );
XOR2X1 XOR2X1_11 ( .A(asr1_dataout_3_), .B(asr2_dataout_3_), .Y(_977_) );
AND2X2 AND2X2_42 ( .A(asr1_dataout_2_), .B(asr2_dataout_2_), .Y(_978_) );
AOI21X1 AOI21X1_65 ( .A(_974_), .B(_975_), .C(_978_), .Y(_979_) );
XOR2X1 XOR2X1_12 ( .A(_979_), .B(_977_), .Y(_980_) );
NOR2X1 NOR2X1_79 ( .A(rst_bF_buf1), .B(_980_), .Y(_963__3_) );
NAND3X1 NAND3X1_248 ( .A(_975_), .B(_977_), .C(_974_), .Y(_981_) );
INVX1 INVX1_214 ( .A(asr1_dataout_3_), .Y(_982_) );
INVX1 INVX1_215 ( .A(asr2_dataout_3_), .Y(_983_) );
NAND2X1 NAND2X1_174 ( .A(_982_), .B(_983_), .Y(_984_) );
NOR2X1 NOR2X1_80 ( .A(_982_), .B(_983_), .Y(_985_) );
AOI21X1 AOI21X1_66 ( .A(_978_), .B(_984_), .C(_985_), .Y(_986_) );
NAND2X1 NAND2X1_175 ( .A(_986_), .B(_981_), .Y(_987_) );
XOR2X1 XOR2X1_13 ( .A(asr1_dataout_4_), .B(asr2_dataout_4_), .Y(_988_) );
OAI21X1 OAI21X1_115 ( .A(_988_), .B(_987_), .C(_966_), .Y(_989_) );
AOI21X1 AOI21X1_67 ( .A(_987_), .B(_988_), .C(_989_), .Y(_963__4_) );
XOR2X1 XOR2X1_14 ( .A(asr1_dataout_5_), .B(asr2_dataout_5_), .Y(_990_) );
NAND2X1 NAND2X1_176 ( .A(_988_), .B(_990_), .Y(_991_) );
AOI21X1 AOI21X1_68 ( .A(_981_), .B(_986_), .C(_991_), .Y(_992_) );
INVX1 INVX1_216 ( .A(asr1_dataout_4_), .Y(_993_) );
INVX1 INVX1_217 ( .A(asr2_dataout_4_), .Y(_994_) );
NAND2X1 NAND2X1_177 ( .A(_988_), .B(_987_), .Y(_995_) );
OAI21X1 OAI21X1_116 ( .A(_993_), .B(_994_), .C(_995_), .Y(_996_) );
NOR2X1 NOR2X1_81 ( .A(_993_), .B(_994_), .Y(_997_) );
AOI21X1 AOI21X1_69 ( .A(_990_), .B(_997_), .C(rst_bF_buf0), .Y(_998_) );
OAI21X1 OAI21X1_117 ( .A(_990_), .B(_996_), .C(_998_), .Y(_999_) );
NOR2X1 NOR2X1_82 ( .A(_992_), .B(_999_), .Y(_963__5_) );
NAND2X1 NAND2X1_178 ( .A(asr1_dataout_5_), .B(asr2_dataout_5_), .Y(_1000_) );
NAND2X1 NAND2X1_179 ( .A(_997_), .B(_990_), .Y(_1001_) );
NAND2X1 NAND2X1_180 ( .A(_1000_), .B(_1001_), .Y(_1002_) );
OR2X2 OR2X2_6 ( .A(_992_), .B(_1002_), .Y(_1003_) );
XOR2X1 XOR2X1_15 ( .A(asr1_dataout_6_), .B(asr2_dataout_6_), .Y(_1004_) );
OAI21X1 OAI21X1_118 ( .A(_1004_), .B(_1003_), .C(_966_), .Y(_1005_) );
AOI21X1 AOI21X1_70 ( .A(_1003_), .B(_1004_), .C(_1005_), .Y(_963__6_) );
NAND2X1 NAND2X1_181 ( .A(asr1_dataout_6_), .B(asr2_dataout_6_), .Y(_1006_) );
OAI21X1 OAI21X1_119 ( .A(_1002_), .B(_992_), .C(_1004_), .Y(_1007_) );
XNOR2X1 XNOR2X1_4 ( .A(asr1_dataout_7_), .B(asr2_dataout_7_), .Y(_1008_) );
AOI21X1 AOI21X1_71 ( .A(_1007_), .B(_1006_), .C(_1008_), .Y(_1009_) );
NAND3X1 NAND3X1_249 ( .A(_1006_), .B(_1008_), .C(_1007_), .Y(_1010_) );
NAND2X1 NAND2X1_182 ( .A(_966_), .B(_1010_), .Y(_1011_) );
NOR2X1 NOR2X1_83 ( .A(_1009_), .B(_1011_), .Y(_963__7_) );
DFFPOSX1 DFFPOSX1_43 ( .CLK(clk_bF_buf6), .D(_963__0_), .Q(sumador_res_0_) );
DFFPOSX1 DFFPOSX1_44 ( .CLK(clk_bF_buf2), .D(_963__1_), .Q(sumador_res_1_) );
DFFPOSX1 DFFPOSX1_45 ( .CLK(clk_bF_buf1), .D(_963__2_), .Q(sumador_res_2_) );
DFFPOSX1 DFFPOSX1_46 ( .CLK(clk_bF_buf0), .D(_963__3_), .Q(sumador_res_3_) );
DFFPOSX1 DFFPOSX1_47 ( .CLK(clk_bF_buf4), .D(_963__4_), .Q(sumador_res_4_) );
DFFPOSX1 DFFPOSX1_48 ( .CLK(clk_bF_buf4), .D(_963__5_), .Q(sumador_res_5_) );
DFFPOSX1 DFFPOSX1_49 ( .CLK(clk_bF_buf3), .D(_963__6_), .Q(sumador_res_6_) );
DFFPOSX1 DFFPOSX1_50 ( .CLK(clk_bF_buf4), .D(_963__7_), .Q(sumador_res_7_) );
BUFX2 BUFX2_79 ( .A(1'b0), .Y(_955__5_) );
BUFX2 BUFX2_80 ( .A(1'b0), .Y(_955__6_) );
BUFX2 BUFX2_81 ( .A(1'b0), .Y(_955__7_) );
BUFX2 BUFX2_82 ( .A(asr1_en_0_), .Y(asr1_rom_15__0_) );
BUFX2 BUFX2_83 ( .A(asr1_en_1_), .Y(asr1_rom_15__1_) );
BUFX2 BUFX2_84 ( .A(asr1_en_2_), .Y(asr1_rom_15__2_) );
BUFX2 BUFX2_85 ( .A(asr1_en_3_), .Y(asr1_rom_15__3_) );
BUFX2 BUFX2_86 ( .A(asr1_en_4_), .Y(asr1_rom_15__4_) );
BUFX2 BUFX2_87 ( .A(asr1_en_5_), .Y(asr1_rom_15__5_) );
BUFX2 BUFX2_88 ( .A(asr1_en_6_), .Y(asr1_rom_15__6_) );
BUFX2 BUFX2_89 ( .A(asr1_en_7_), .Y(asr1_rom_15__7_) );
BUFX2 BUFX2_90 ( .A(asr2_en_0_), .Y(asr2_rom_15__0_) );
BUFX2 BUFX2_91 ( .A(asr2_en_1_), .Y(asr2_rom_15__1_) );
BUFX2 BUFX2_92 ( .A(asr2_en_2_), .Y(asr2_rom_15__2_) );
BUFX2 BUFX2_93 ( .A(asr2_en_3_), .Y(asr2_rom_15__3_) );
BUFX2 BUFX2_94 ( .A(asr2_en_4_), .Y(asr2_rom_15__4_) );
BUFX2 BUFX2_95 ( .A(asr2_en_5_), .Y(asr2_rom_15__5_) );
BUFX2 BUFX2_96 ( .A(asr2_en_6_), .Y(asr2_rom_15__6_) );
BUFX2 BUFX2_97 ( .A(asr2_en_7_), .Y(asr2_rom_15__7_) );
BUFX2 BUFX2_98 ( .A(1'b0), .Y(rom1_data_5_) );
BUFX2 BUFX2_99 ( .A(1'b0), .Y(rom1_data_6_) );
BUFX2 BUFX2_100 ( .A(1'b0), .Y(rom1_data_7_) );
FILL FILL_0_DFFSR_274 ( );
FILL FILL_1_DFFSR_274 ( );
FILL FILL_2_DFFSR_274 ( );
FILL FILL_3_DFFSR_274 ( );
FILL FILL_4_DFFSR_274 ( );
FILL FILL_5_DFFSR_274 ( );
FILL FILL_6_DFFSR_274 ( );
FILL FILL_7_DFFSR_274 ( );
FILL FILL_8_DFFSR_274 ( );
FILL FILL_9_DFFSR_274 ( );
FILL FILL_10_DFFSR_274 ( );
FILL FILL_11_DFFSR_274 ( );
FILL FILL_12_DFFSR_274 ( );
FILL FILL_13_DFFSR_274 ( );
FILL FILL_14_DFFSR_274 ( );
FILL FILL_15_DFFSR_274 ( );
FILL FILL_16_DFFSR_274 ( );
FILL FILL_17_DFFSR_274 ( );
FILL FILL_18_DFFSR_274 ( );
FILL FILL_19_DFFSR_274 ( );
FILL FILL_20_DFFSR_274 ( );
FILL FILL_21_DFFSR_274 ( );
FILL FILL_22_DFFSR_274 ( );
FILL FILL_23_DFFSR_274 ( );
FILL FILL_24_DFFSR_274 ( );
FILL FILL_25_DFFSR_274 ( );
FILL FILL_26_DFFSR_274 ( );
FILL FILL_27_DFFSR_274 ( );
FILL FILL_28_DFFSR_274 ( );
FILL FILL_29_DFFSR_274 ( );
FILL FILL_30_DFFSR_274 ( );
FILL FILL_31_DFFSR_274 ( );
FILL FILL_32_DFFSR_274 ( );
FILL FILL_33_DFFSR_274 ( );
FILL FILL_34_DFFSR_274 ( );
FILL FILL_35_DFFSR_274 ( );
FILL FILL_36_DFFSR_274 ( );
FILL FILL_37_DFFSR_274 ( );
FILL FILL_38_DFFSR_274 ( );
FILL FILL_39_DFFSR_274 ( );
FILL FILL_40_DFFSR_274 ( );
FILL FILL_41_DFFSR_274 ( );
FILL FILL_42_DFFSR_274 ( );
FILL FILL_43_DFFSR_274 ( );
FILL FILL_44_DFFSR_274 ( );
FILL FILL_45_DFFSR_274 ( );
FILL FILL_46_DFFSR_274 ( );
FILL FILL_47_DFFSR_274 ( );
FILL FILL_48_DFFSR_274 ( );
FILL FILL_49_DFFSR_274 ( );
FILL FILL_50_DFFSR_274 ( );
FILL FILL_0_NAND2X1_136 ( );
FILL FILL_1_NAND2X1_136 ( );
FILL FILL_2_NAND2X1_136 ( );
FILL FILL_3_NAND2X1_136 ( );
FILL FILL_4_NAND2X1_136 ( );
FILL FILL_5_NAND2X1_136 ( );
FILL FILL_6_NAND2X1_136 ( );
FILL FILL_0_OAI21X1_105 ( );
FILL FILL_1_OAI21X1_105 ( );
FILL FILL_2_OAI21X1_105 ( );
FILL FILL_3_OAI21X1_105 ( );
FILL FILL_4_OAI21X1_105 ( );
FILL FILL_5_OAI21X1_105 ( );
FILL FILL_6_OAI21X1_105 ( );
FILL FILL_7_OAI21X1_105 ( );
FILL FILL_8_OAI21X1_105 ( );
FILL FILL_0_INVX1_194 ( );
FILL FILL_1_INVX1_194 ( );
FILL FILL_2_INVX1_194 ( );
FILL FILL_3_INVX1_194 ( );
FILL FILL_0_OAI21X1_97 ( );
FILL FILL_1_OAI21X1_97 ( );
FILL FILL_2_OAI21X1_97 ( );
FILL FILL_3_OAI21X1_97 ( );
FILL FILL_4_OAI21X1_97 ( );
FILL FILL_5_OAI21X1_97 ( );
FILL FILL_6_OAI21X1_97 ( );
FILL FILL_7_OAI21X1_97 ( );
FILL FILL_8_OAI21X1_97 ( );
FILL FILL_9_OAI21X1_97 ( );
FILL FILL_0_NAND2X1_128 ( );
FILL FILL_1_NAND2X1_128 ( );
FILL FILL_2_NAND2X1_128 ( );
FILL FILL_3_NAND2X1_128 ( );
FILL FILL_4_NAND2X1_128 ( );
FILL FILL_5_NAND2X1_128 ( );
FILL FILL_6_NAND2X1_128 ( );
FILL FILL_0_INVX1_203 ( );
FILL FILL_1_INVX1_203 ( );
FILL FILL_2_INVX1_203 ( );
FILL FILL_3_INVX1_203 ( );
FILL FILL_4_INVX1_203 ( );
FILL FILL_0_BUFX2_75 ( );
FILL FILL_1_BUFX2_75 ( );
FILL FILL_2_BUFX2_75 ( );
FILL FILL_3_BUFX2_75 ( );
FILL FILL_4_BUFX2_75 ( );
FILL FILL_5_BUFX2_75 ( );
FILL FILL_6_BUFX2_75 ( );
FILL FILL_0_DFFPOSX1_29 ( );
FILL FILL_1_DFFPOSX1_29 ( );
FILL FILL_2_DFFPOSX1_29 ( );
FILL FILL_3_DFFPOSX1_29 ( );
FILL FILL_4_DFFPOSX1_29 ( );
FILL FILL_5_DFFPOSX1_29 ( );
FILL FILL_6_DFFPOSX1_29 ( );
FILL FILL_7_DFFPOSX1_29 ( );
FILL FILL_8_DFFPOSX1_29 ( );
FILL FILL_9_DFFPOSX1_29 ( );
FILL FILL_10_DFFPOSX1_29 ( );
FILL FILL_11_DFFPOSX1_29 ( );
FILL FILL_12_DFFPOSX1_29 ( );
FILL FILL_13_DFFPOSX1_29 ( );
FILL FILL_14_DFFPOSX1_29 ( );
FILL FILL_15_DFFPOSX1_29 ( );
FILL FILL_16_DFFPOSX1_29 ( );
FILL FILL_17_DFFPOSX1_29 ( );
FILL FILL_18_DFFPOSX1_29 ( );
FILL FILL_19_DFFPOSX1_29 ( );
FILL FILL_20_DFFPOSX1_29 ( );
FILL FILL_21_DFFPOSX1_29 ( );
FILL FILL_22_DFFPOSX1_29 ( );
FILL FILL_23_DFFPOSX1_29 ( );
FILL FILL_24_DFFPOSX1_29 ( );
FILL FILL_25_DFFPOSX1_29 ( );
FILL FILL_26_DFFPOSX1_29 ( );
FILL FILL_27_DFFPOSX1_29 ( );
FILL FILL_0_DFFSR_276 ( );
FILL FILL_1_DFFSR_276 ( );
FILL FILL_2_DFFSR_276 ( );
FILL FILL_3_DFFSR_276 ( );
FILL FILL_4_DFFSR_276 ( );
FILL FILL_5_DFFSR_276 ( );
FILL FILL_6_DFFSR_276 ( );
FILL FILL_7_DFFSR_276 ( );
FILL FILL_8_DFFSR_276 ( );
FILL FILL_9_DFFSR_276 ( );
FILL FILL_10_DFFSR_276 ( );
FILL FILL_11_DFFSR_276 ( );
FILL FILL_12_DFFSR_276 ( );
FILL FILL_13_DFFSR_276 ( );
FILL FILL_14_DFFSR_276 ( );
FILL FILL_15_DFFSR_276 ( );
FILL FILL_16_DFFSR_276 ( );
FILL FILL_17_DFFSR_276 ( );
FILL FILL_18_DFFSR_276 ( );
FILL FILL_19_DFFSR_276 ( );
FILL FILL_20_DFFSR_276 ( );
FILL FILL_21_DFFSR_276 ( );
FILL FILL_22_DFFSR_276 ( );
FILL FILL_23_DFFSR_276 ( );
FILL FILL_24_DFFSR_276 ( );
FILL FILL_25_DFFSR_276 ( );
FILL FILL_26_DFFSR_276 ( );
FILL FILL_27_DFFSR_276 ( );
FILL FILL_28_DFFSR_276 ( );
FILL FILL_29_DFFSR_276 ( );
FILL FILL_30_DFFSR_276 ( );
FILL FILL_31_DFFSR_276 ( );
FILL FILL_32_DFFSR_276 ( );
FILL FILL_33_DFFSR_276 ( );
FILL FILL_34_DFFSR_276 ( );
FILL FILL_35_DFFSR_276 ( );
FILL FILL_36_DFFSR_276 ( );
FILL FILL_37_DFFSR_276 ( );
FILL FILL_38_DFFSR_276 ( );
FILL FILL_39_DFFSR_276 ( );
FILL FILL_40_DFFSR_276 ( );
FILL FILL_41_DFFSR_276 ( );
FILL FILL_42_DFFSR_276 ( );
FILL FILL_43_DFFSR_276 ( );
FILL FILL_44_DFFSR_276 ( );
FILL FILL_45_DFFSR_276 ( );
FILL FILL_46_DFFSR_276 ( );
FILL FILL_47_DFFSR_276 ( );
FILL FILL_48_DFFSR_276 ( );
FILL FILL_49_DFFSR_276 ( );
FILL FILL_50_DFFSR_276 ( );
FILL FILL_0_BUFX2_74 ( );
FILL FILL_1_BUFX2_74 ( );
FILL FILL_2_BUFX2_74 ( );
FILL FILL_3_BUFX2_74 ( );
FILL FILL_4_BUFX2_74 ( );
FILL FILL_5_BUFX2_74 ( );
FILL FILL_6_BUFX2_74 ( );
FILL FILL_0_DFFSR_214 ( );
FILL FILL_1_DFFSR_214 ( );
FILL FILL_2_DFFSR_214 ( );
FILL FILL_3_DFFSR_214 ( );
FILL FILL_4_DFFSR_214 ( );
FILL FILL_5_DFFSR_214 ( );
FILL FILL_6_DFFSR_214 ( );
FILL FILL_7_DFFSR_214 ( );
FILL FILL_8_DFFSR_214 ( );
FILL FILL_9_DFFSR_214 ( );
FILL FILL_10_DFFSR_214 ( );
FILL FILL_11_DFFSR_214 ( );
FILL FILL_12_DFFSR_214 ( );
FILL FILL_13_DFFSR_214 ( );
FILL FILL_14_DFFSR_214 ( );
FILL FILL_15_DFFSR_214 ( );
FILL FILL_16_DFFSR_214 ( );
FILL FILL_17_DFFSR_214 ( );
FILL FILL_18_DFFSR_214 ( );
FILL FILL_19_DFFSR_214 ( );
FILL FILL_20_DFFSR_214 ( );
FILL FILL_21_DFFSR_214 ( );
FILL FILL_22_DFFSR_214 ( );
FILL FILL_23_DFFSR_214 ( );
FILL FILL_24_DFFSR_214 ( );
FILL FILL_25_DFFSR_214 ( );
FILL FILL_26_DFFSR_214 ( );
FILL FILL_27_DFFSR_214 ( );
FILL FILL_28_DFFSR_214 ( );
FILL FILL_29_DFFSR_214 ( );
FILL FILL_30_DFFSR_214 ( );
FILL FILL_31_DFFSR_214 ( );
FILL FILL_32_DFFSR_214 ( );
FILL FILL_33_DFFSR_214 ( );
FILL FILL_34_DFFSR_214 ( );
FILL FILL_35_DFFSR_214 ( );
FILL FILL_36_DFFSR_214 ( );
FILL FILL_37_DFFSR_214 ( );
FILL FILL_38_DFFSR_214 ( );
FILL FILL_39_DFFSR_214 ( );
FILL FILL_40_DFFSR_214 ( );
FILL FILL_41_DFFSR_214 ( );
FILL FILL_42_DFFSR_214 ( );
FILL FILL_43_DFFSR_214 ( );
FILL FILL_44_DFFSR_214 ( );
FILL FILL_45_DFFSR_214 ( );
FILL FILL_46_DFFSR_214 ( );
FILL FILL_47_DFFSR_214 ( );
FILL FILL_48_DFFSR_214 ( );
FILL FILL_49_DFFSR_214 ( );
FILL FILL_50_DFFSR_214 ( );
FILL FILL_51_DFFSR_214 ( );
FILL FILL_0_DFFSR_238 ( );
FILL FILL_1_DFFSR_238 ( );
FILL FILL_2_DFFSR_238 ( );
FILL FILL_3_DFFSR_238 ( );
FILL FILL_4_DFFSR_238 ( );
FILL FILL_5_DFFSR_238 ( );
FILL FILL_6_DFFSR_238 ( );
FILL FILL_7_DFFSR_238 ( );
FILL FILL_8_DFFSR_238 ( );
FILL FILL_9_DFFSR_238 ( );
FILL FILL_10_DFFSR_238 ( );
FILL FILL_11_DFFSR_238 ( );
FILL FILL_12_DFFSR_238 ( );
FILL FILL_13_DFFSR_238 ( );
FILL FILL_14_DFFSR_238 ( );
FILL FILL_15_DFFSR_238 ( );
FILL FILL_16_DFFSR_238 ( );
FILL FILL_17_DFFSR_238 ( );
FILL FILL_18_DFFSR_238 ( );
FILL FILL_19_DFFSR_238 ( );
FILL FILL_20_DFFSR_238 ( );
FILL FILL_21_DFFSR_238 ( );
FILL FILL_22_DFFSR_238 ( );
FILL FILL_23_DFFSR_238 ( );
FILL FILL_24_DFFSR_238 ( );
FILL FILL_25_DFFSR_238 ( );
FILL FILL_26_DFFSR_238 ( );
FILL FILL_27_DFFSR_238 ( );
FILL FILL_28_DFFSR_238 ( );
FILL FILL_29_DFFSR_238 ( );
FILL FILL_30_DFFSR_238 ( );
FILL FILL_31_DFFSR_238 ( );
FILL FILL_32_DFFSR_238 ( );
FILL FILL_33_DFFSR_238 ( );
FILL FILL_34_DFFSR_238 ( );
FILL FILL_35_DFFSR_238 ( );
FILL FILL_36_DFFSR_238 ( );
FILL FILL_37_DFFSR_238 ( );
FILL FILL_38_DFFSR_238 ( );
FILL FILL_39_DFFSR_238 ( );
FILL FILL_40_DFFSR_238 ( );
FILL FILL_41_DFFSR_238 ( );
FILL FILL_42_DFFSR_238 ( );
FILL FILL_43_DFFSR_238 ( );
FILL FILL_44_DFFSR_238 ( );
FILL FILL_45_DFFSR_238 ( );
FILL FILL_46_DFFSR_238 ( );
FILL FILL_47_DFFSR_238 ( );
FILL FILL_48_DFFSR_238 ( );
FILL FILL_49_DFFSR_238 ( );
FILL FILL_50_DFFSR_238 ( );
FILL FILL_0_DFFSR_249 ( );
FILL FILL_1_DFFSR_249 ( );
FILL FILL_2_DFFSR_249 ( );
FILL FILL_3_DFFSR_249 ( );
FILL FILL_4_DFFSR_249 ( );
FILL FILL_5_DFFSR_249 ( );
FILL FILL_6_DFFSR_249 ( );
FILL FILL_7_DFFSR_249 ( );
FILL FILL_8_DFFSR_249 ( );
FILL FILL_9_DFFSR_249 ( );
FILL FILL_10_DFFSR_249 ( );
FILL FILL_11_DFFSR_249 ( );
FILL FILL_12_DFFSR_249 ( );
FILL FILL_13_DFFSR_249 ( );
FILL FILL_14_DFFSR_249 ( );
FILL FILL_15_DFFSR_249 ( );
FILL FILL_16_DFFSR_249 ( );
FILL FILL_17_DFFSR_249 ( );
FILL FILL_18_DFFSR_249 ( );
FILL FILL_19_DFFSR_249 ( );
FILL FILL_20_DFFSR_249 ( );
FILL FILL_21_DFFSR_249 ( );
FILL FILL_22_DFFSR_249 ( );
FILL FILL_23_DFFSR_249 ( );
FILL FILL_24_DFFSR_249 ( );
FILL FILL_25_DFFSR_249 ( );
FILL FILL_26_DFFSR_249 ( );
FILL FILL_27_DFFSR_249 ( );
FILL FILL_28_DFFSR_249 ( );
FILL FILL_29_DFFSR_249 ( );
FILL FILL_30_DFFSR_249 ( );
FILL FILL_31_DFFSR_249 ( );
FILL FILL_32_DFFSR_249 ( );
FILL FILL_33_DFFSR_249 ( );
FILL FILL_34_DFFSR_249 ( );
FILL FILL_35_DFFSR_249 ( );
FILL FILL_36_DFFSR_249 ( );
FILL FILL_37_DFFSR_249 ( );
FILL FILL_38_DFFSR_249 ( );
FILL FILL_39_DFFSR_249 ( );
FILL FILL_40_DFFSR_249 ( );
FILL FILL_41_DFFSR_249 ( );
FILL FILL_42_DFFSR_249 ( );
FILL FILL_43_DFFSR_249 ( );
FILL FILL_44_DFFSR_249 ( );
FILL FILL_45_DFFSR_249 ( );
FILL FILL_46_DFFSR_249 ( );
FILL FILL_47_DFFSR_249 ( );
FILL FILL_48_DFFSR_249 ( );
FILL FILL_49_DFFSR_249 ( );
FILL FILL_50_DFFSR_249 ( );
FILL FILL_0_CLKBUF1_2 ( );
FILL FILL_1_CLKBUF1_2 ( );
FILL FILL_2_CLKBUF1_2 ( );
FILL FILL_3_CLKBUF1_2 ( );
FILL FILL_4_CLKBUF1_2 ( );
FILL FILL_5_CLKBUF1_2 ( );
FILL FILL_6_CLKBUF1_2 ( );
FILL FILL_7_CLKBUF1_2 ( );
FILL FILL_8_CLKBUF1_2 ( );
FILL FILL_9_CLKBUF1_2 ( );
FILL FILL_10_CLKBUF1_2 ( );
FILL FILL_11_CLKBUF1_2 ( );
FILL FILL_12_CLKBUF1_2 ( );
FILL FILL_13_CLKBUF1_2 ( );
FILL FILL_14_CLKBUF1_2 ( );
FILL FILL_15_CLKBUF1_2 ( );
FILL FILL_16_CLKBUF1_2 ( );
FILL FILL_17_CLKBUF1_2 ( );
FILL FILL_18_CLKBUF1_2 ( );
FILL FILL_19_CLKBUF1_2 ( );
FILL FILL_20_CLKBUF1_2 ( );
FILL FILL_0_DFFSR_209 ( );
FILL FILL_1_DFFSR_209 ( );
FILL FILL_2_DFFSR_209 ( );
FILL FILL_3_DFFSR_209 ( );
FILL FILL_4_DFFSR_209 ( );
FILL FILL_5_DFFSR_209 ( );
FILL FILL_6_DFFSR_209 ( );
FILL FILL_7_DFFSR_209 ( );
FILL FILL_8_DFFSR_209 ( );
FILL FILL_9_DFFSR_209 ( );
FILL FILL_10_DFFSR_209 ( );
FILL FILL_11_DFFSR_209 ( );
FILL FILL_12_DFFSR_209 ( );
FILL FILL_13_DFFSR_209 ( );
FILL FILL_14_DFFSR_209 ( );
FILL FILL_15_DFFSR_209 ( );
FILL FILL_16_DFFSR_209 ( );
FILL FILL_17_DFFSR_209 ( );
FILL FILL_18_DFFSR_209 ( );
FILL FILL_19_DFFSR_209 ( );
FILL FILL_20_DFFSR_209 ( );
FILL FILL_21_DFFSR_209 ( );
FILL FILL_22_DFFSR_209 ( );
FILL FILL_23_DFFSR_209 ( );
FILL FILL_24_DFFSR_209 ( );
FILL FILL_25_DFFSR_209 ( );
FILL FILL_26_DFFSR_209 ( );
FILL FILL_27_DFFSR_209 ( );
FILL FILL_28_DFFSR_209 ( );
FILL FILL_29_DFFSR_209 ( );
FILL FILL_30_DFFSR_209 ( );
FILL FILL_31_DFFSR_209 ( );
FILL FILL_32_DFFSR_209 ( );
FILL FILL_33_DFFSR_209 ( );
FILL FILL_34_DFFSR_209 ( );
FILL FILL_35_DFFSR_209 ( );
FILL FILL_36_DFFSR_209 ( );
FILL FILL_37_DFFSR_209 ( );
FILL FILL_38_DFFSR_209 ( );
FILL FILL_39_DFFSR_209 ( );
FILL FILL_40_DFFSR_209 ( );
FILL FILL_41_DFFSR_209 ( );
FILL FILL_42_DFFSR_209 ( );
FILL FILL_43_DFFSR_209 ( );
FILL FILL_44_DFFSR_209 ( );
FILL FILL_45_DFFSR_209 ( );
FILL FILL_46_DFFSR_209 ( );
FILL FILL_47_DFFSR_209 ( );
FILL FILL_48_DFFSR_209 ( );
FILL FILL_49_DFFSR_209 ( );
FILL FILL_50_DFFSR_209 ( );
FILL FILL_0_OAI22X1_45 ( );
FILL FILL_1_OAI22X1_45 ( );
FILL FILL_2_OAI22X1_45 ( );
FILL FILL_3_OAI22X1_45 ( );
FILL FILL_4_OAI22X1_45 ( );
FILL FILL_5_OAI22X1_45 ( );
FILL FILL_6_OAI22X1_45 ( );
FILL FILL_7_OAI22X1_45 ( );
FILL FILL_8_OAI22X1_45 ( );
FILL FILL_9_OAI22X1_45 ( );
FILL FILL_10_OAI22X1_45 ( );
FILL FILL_11_OAI22X1_45 ( );
FILL FILL_0_DFFSR_149 ( );
FILL FILL_1_DFFSR_149 ( );
FILL FILL_2_DFFSR_149 ( );
FILL FILL_3_DFFSR_149 ( );
FILL FILL_4_DFFSR_149 ( );
FILL FILL_5_DFFSR_149 ( );
FILL FILL_6_DFFSR_149 ( );
FILL FILL_7_DFFSR_149 ( );
FILL FILL_8_DFFSR_149 ( );
FILL FILL_9_DFFSR_149 ( );
FILL FILL_10_DFFSR_149 ( );
FILL FILL_11_DFFSR_149 ( );
FILL FILL_12_DFFSR_149 ( );
FILL FILL_13_DFFSR_149 ( );
FILL FILL_14_DFFSR_149 ( );
FILL FILL_15_DFFSR_149 ( );
FILL FILL_16_DFFSR_149 ( );
FILL FILL_17_DFFSR_149 ( );
FILL FILL_18_DFFSR_149 ( );
FILL FILL_19_DFFSR_149 ( );
FILL FILL_20_DFFSR_149 ( );
FILL FILL_21_DFFSR_149 ( );
FILL FILL_22_DFFSR_149 ( );
FILL FILL_23_DFFSR_149 ( );
FILL FILL_24_DFFSR_149 ( );
FILL FILL_25_DFFSR_149 ( );
FILL FILL_26_DFFSR_149 ( );
FILL FILL_27_DFFSR_149 ( );
FILL FILL_28_DFFSR_149 ( );
FILL FILL_29_DFFSR_149 ( );
FILL FILL_30_DFFSR_149 ( );
FILL FILL_31_DFFSR_149 ( );
FILL FILL_32_DFFSR_149 ( );
FILL FILL_33_DFFSR_149 ( );
FILL FILL_34_DFFSR_149 ( );
FILL FILL_35_DFFSR_149 ( );
FILL FILL_36_DFFSR_149 ( );
FILL FILL_37_DFFSR_149 ( );
FILL FILL_38_DFFSR_149 ( );
FILL FILL_39_DFFSR_149 ( );
FILL FILL_40_DFFSR_149 ( );
FILL FILL_41_DFFSR_149 ( );
FILL FILL_42_DFFSR_149 ( );
FILL FILL_43_DFFSR_149 ( );
FILL FILL_44_DFFSR_149 ( );
FILL FILL_45_DFFSR_149 ( );
FILL FILL_46_DFFSR_149 ( );
FILL FILL_47_DFFSR_149 ( );
FILL FILL_48_DFFSR_149 ( );
FILL FILL_49_DFFSR_149 ( );
FILL FILL_50_DFFSR_149 ( );
FILL FILL_51_DFFSR_149 ( );
FILL FILL_0_NAND2X1_133 ( );
FILL FILL_1_NAND2X1_133 ( );
FILL FILL_2_NAND2X1_133 ( );
FILL FILL_3_NAND2X1_133 ( );
FILL FILL_4_NAND2X1_133 ( );
FILL FILL_5_NAND2X1_133 ( );
FILL FILL_6_NAND2X1_133 ( );
FILL FILL_0_OAI21X1_102 ( );
FILL FILL_1_OAI21X1_102 ( );
FILL FILL_2_OAI21X1_102 ( );
FILL FILL_3_OAI21X1_102 ( );
FILL FILL_4_OAI21X1_102 ( );
FILL FILL_5_OAI21X1_102 ( );
FILL FILL_6_OAI21X1_102 ( );
FILL FILL_7_OAI21X1_102 ( );
FILL FILL_8_OAI21X1_102 ( );
FILL FILL_0_INVX1_200 ( );
FILL FILL_1_INVX1_200 ( );
FILL FILL_2_INVX1_200 ( );
FILL FILL_3_INVX1_200 ( );
FILL FILL_4_INVX1_200 ( );
FILL FILL_0_BUFX2_72 ( );
FILL FILL_1_BUFX2_72 ( );
FILL FILL_2_BUFX2_72 ( );
FILL FILL_3_BUFX2_72 ( );
FILL FILL_4_BUFX2_72 ( );
FILL FILL_5_BUFX2_72 ( );
FILL FILL_6_BUFX2_72 ( );
FILL FILL_0_DFFPOSX1_15 ( );
FILL FILL_1_DFFPOSX1_15 ( );
FILL FILL_2_DFFPOSX1_15 ( );
FILL FILL_3_DFFPOSX1_15 ( );
FILL FILL_4_DFFPOSX1_15 ( );
FILL FILL_5_DFFPOSX1_15 ( );
FILL FILL_6_DFFPOSX1_15 ( );
FILL FILL_7_DFFPOSX1_15 ( );
FILL FILL_8_DFFPOSX1_15 ( );
FILL FILL_9_DFFPOSX1_15 ( );
FILL FILL_10_DFFPOSX1_15 ( );
FILL FILL_11_DFFPOSX1_15 ( );
FILL FILL_12_DFFPOSX1_15 ( );
FILL FILL_13_DFFPOSX1_15 ( );
FILL FILL_14_DFFPOSX1_15 ( );
FILL FILL_15_DFFPOSX1_15 ( );
FILL FILL_16_DFFPOSX1_15 ( );
FILL FILL_17_DFFPOSX1_15 ( );
FILL FILL_18_DFFPOSX1_15 ( );
FILL FILL_19_DFFPOSX1_15 ( );
FILL FILL_20_DFFPOSX1_15 ( );
FILL FILL_21_DFFPOSX1_15 ( );
FILL FILL_22_DFFPOSX1_15 ( );
FILL FILL_23_DFFPOSX1_15 ( );
FILL FILL_24_DFFPOSX1_15 ( );
FILL FILL_25_DFFPOSX1_15 ( );
FILL FILL_26_DFFPOSX1_15 ( );
FILL FILL_27_DFFPOSX1_15 ( );
FILL FILL_0_DFFSR_277 ( );
FILL FILL_1_DFFSR_277 ( );
FILL FILL_2_DFFSR_277 ( );
FILL FILL_3_DFFSR_277 ( );
FILL FILL_4_DFFSR_277 ( );
FILL FILL_5_DFFSR_277 ( );
FILL FILL_6_DFFSR_277 ( );
FILL FILL_7_DFFSR_277 ( );
FILL FILL_8_DFFSR_277 ( );
FILL FILL_9_DFFSR_277 ( );
FILL FILL_10_DFFSR_277 ( );
FILL FILL_11_DFFSR_277 ( );
FILL FILL_12_DFFSR_277 ( );
FILL FILL_13_DFFSR_277 ( );
FILL FILL_14_DFFSR_277 ( );
FILL FILL_15_DFFSR_277 ( );
FILL FILL_16_DFFSR_277 ( );
FILL FILL_17_DFFSR_277 ( );
FILL FILL_18_DFFSR_277 ( );
FILL FILL_19_DFFSR_277 ( );
FILL FILL_20_DFFSR_277 ( );
FILL FILL_21_DFFSR_277 ( );
FILL FILL_22_DFFSR_277 ( );
FILL FILL_23_DFFSR_277 ( );
FILL FILL_24_DFFSR_277 ( );
FILL FILL_25_DFFSR_277 ( );
FILL FILL_26_DFFSR_277 ( );
FILL FILL_27_DFFSR_277 ( );
FILL FILL_28_DFFSR_277 ( );
FILL FILL_29_DFFSR_277 ( );
FILL FILL_30_DFFSR_277 ( );
FILL FILL_31_DFFSR_277 ( );
FILL FILL_32_DFFSR_277 ( );
FILL FILL_33_DFFSR_277 ( );
FILL FILL_34_DFFSR_277 ( );
FILL FILL_35_DFFSR_277 ( );
FILL FILL_36_DFFSR_277 ( );
FILL FILL_37_DFFSR_277 ( );
FILL FILL_38_DFFSR_277 ( );
FILL FILL_39_DFFSR_277 ( );
FILL FILL_40_DFFSR_277 ( );
FILL FILL_41_DFFSR_277 ( );
FILL FILL_42_DFFSR_277 ( );
FILL FILL_43_DFFSR_277 ( );
FILL FILL_44_DFFSR_277 ( );
FILL FILL_45_DFFSR_277 ( );
FILL FILL_46_DFFSR_277 ( );
FILL FILL_47_DFFSR_277 ( );
FILL FILL_48_DFFSR_277 ( );
FILL FILL_49_DFFSR_277 ( );
FILL FILL_50_DFFSR_277 ( );
FILL FILL_0_NAND2X1_161 ( );
FILL FILL_1_NAND2X1_161 ( );
FILL FILL_2_NAND2X1_161 ( );
FILL FILL_3_NAND2X1_161 ( );
FILL FILL_4_NAND2X1_161 ( );
FILL FILL_5_NAND2X1_161 ( );
FILL FILL_6_NAND2X1_161 ( );
FILL FILL_0_NAND2X1_162 ( );
FILL FILL_1_NAND2X1_162 ( );
FILL FILL_2_NAND2X1_162 ( );
FILL FILL_3_NAND2X1_162 ( );
FILL FILL_4_NAND2X1_162 ( );
FILL FILL_5_NAND2X1_162 ( );
FILL FILL_6_NAND2X1_162 ( );
FILL FILL_0_DFFPOSX1_37 ( );
FILL FILL_1_DFFPOSX1_37 ( );
FILL FILL_2_DFFPOSX1_37 ( );
FILL FILL_3_DFFPOSX1_37 ( );
FILL FILL_4_DFFPOSX1_37 ( );
FILL FILL_5_DFFPOSX1_37 ( );
FILL FILL_6_DFFPOSX1_37 ( );
FILL FILL_7_DFFPOSX1_37 ( );
FILL FILL_8_DFFPOSX1_37 ( );
FILL FILL_9_DFFPOSX1_37 ( );
FILL FILL_10_DFFPOSX1_37 ( );
FILL FILL_11_DFFPOSX1_37 ( );
FILL FILL_12_DFFPOSX1_37 ( );
FILL FILL_13_DFFPOSX1_37 ( );
FILL FILL_14_DFFPOSX1_37 ( );
FILL FILL_15_DFFPOSX1_37 ( );
FILL FILL_16_DFFPOSX1_37 ( );
FILL FILL_17_DFFPOSX1_37 ( );
FILL FILL_18_DFFPOSX1_37 ( );
FILL FILL_19_DFFPOSX1_37 ( );
FILL FILL_20_DFFPOSX1_37 ( );
FILL FILL_21_DFFPOSX1_37 ( );
FILL FILL_22_DFFPOSX1_37 ( );
FILL FILL_23_DFFPOSX1_37 ( );
FILL FILL_24_DFFPOSX1_37 ( );
FILL FILL_25_DFFPOSX1_37 ( );
FILL FILL_26_DFFPOSX1_37 ( );
FILL FILL_27_DFFPOSX1_37 ( );
FILL FILL_0_INVX1_202 ( );
FILL FILL_1_INVX1_202 ( );
FILL FILL_2_INVX1_202 ( );
FILL FILL_3_INVX1_202 ( );
FILL FILL_4_INVX1_202 ( );
FILL FILL_0_DFFPOSX1_28 ( );
FILL FILL_1_DFFPOSX1_28 ( );
FILL FILL_2_DFFPOSX1_28 ( );
FILL FILL_3_DFFPOSX1_28 ( );
FILL FILL_4_DFFPOSX1_28 ( );
FILL FILL_5_DFFPOSX1_28 ( );
FILL FILL_6_DFFPOSX1_28 ( );
FILL FILL_7_DFFPOSX1_28 ( );
FILL FILL_8_DFFPOSX1_28 ( );
FILL FILL_9_DFFPOSX1_28 ( );
FILL FILL_10_DFFPOSX1_28 ( );
FILL FILL_11_DFFPOSX1_28 ( );
FILL FILL_12_DFFPOSX1_28 ( );
FILL FILL_13_DFFPOSX1_28 ( );
FILL FILL_14_DFFPOSX1_28 ( );
FILL FILL_15_DFFPOSX1_28 ( );
FILL FILL_16_DFFPOSX1_28 ( );
FILL FILL_17_DFFPOSX1_28 ( );
FILL FILL_18_DFFPOSX1_28 ( );
FILL FILL_19_DFFPOSX1_28 ( );
FILL FILL_20_DFFPOSX1_28 ( );
FILL FILL_21_DFFPOSX1_28 ( );
FILL FILL_22_DFFPOSX1_28 ( );
FILL FILL_23_DFFPOSX1_28 ( );
FILL FILL_24_DFFPOSX1_28 ( );
FILL FILL_25_DFFPOSX1_28 ( );
FILL FILL_26_DFFPOSX1_28 ( );
FILL FILL_27_DFFPOSX1_28 ( );
FILL FILL_0_CLKBUF1_31 ( );
FILL FILL_1_CLKBUF1_31 ( );
FILL FILL_2_CLKBUF1_31 ( );
FILL FILL_3_CLKBUF1_31 ( );
FILL FILL_4_CLKBUF1_31 ( );
FILL FILL_5_CLKBUF1_31 ( );
FILL FILL_6_CLKBUF1_31 ( );
FILL FILL_7_CLKBUF1_31 ( );
FILL FILL_8_CLKBUF1_31 ( );
FILL FILL_9_CLKBUF1_31 ( );
FILL FILL_10_CLKBUF1_31 ( );
FILL FILL_11_CLKBUF1_31 ( );
FILL FILL_12_CLKBUF1_31 ( );
FILL FILL_13_CLKBUF1_31 ( );
FILL FILL_14_CLKBUF1_31 ( );
FILL FILL_15_CLKBUF1_31 ( );
FILL FILL_16_CLKBUF1_31 ( );
FILL FILL_17_CLKBUF1_31 ( );
FILL FILL_18_CLKBUF1_31 ( );
FILL FILL_19_CLKBUF1_31 ( );
FILL FILL_20_CLKBUF1_31 ( );
FILL FILL_0_DFFSR_222 ( );
FILL FILL_1_DFFSR_222 ( );
FILL FILL_2_DFFSR_222 ( );
FILL FILL_3_DFFSR_222 ( );
FILL FILL_4_DFFSR_222 ( );
FILL FILL_5_DFFSR_222 ( );
FILL FILL_6_DFFSR_222 ( );
FILL FILL_7_DFFSR_222 ( );
FILL FILL_8_DFFSR_222 ( );
FILL FILL_9_DFFSR_222 ( );
FILL FILL_10_DFFSR_222 ( );
FILL FILL_11_DFFSR_222 ( );
FILL FILL_12_DFFSR_222 ( );
FILL FILL_13_DFFSR_222 ( );
FILL FILL_14_DFFSR_222 ( );
FILL FILL_15_DFFSR_222 ( );
FILL FILL_16_DFFSR_222 ( );
FILL FILL_17_DFFSR_222 ( );
FILL FILL_18_DFFSR_222 ( );
FILL FILL_19_DFFSR_222 ( );
FILL FILL_20_DFFSR_222 ( );
FILL FILL_21_DFFSR_222 ( );
FILL FILL_22_DFFSR_222 ( );
FILL FILL_23_DFFSR_222 ( );
FILL FILL_24_DFFSR_222 ( );
FILL FILL_25_DFFSR_222 ( );
FILL FILL_26_DFFSR_222 ( );
FILL FILL_27_DFFSR_222 ( );
FILL FILL_28_DFFSR_222 ( );
FILL FILL_29_DFFSR_222 ( );
FILL FILL_30_DFFSR_222 ( );
FILL FILL_31_DFFSR_222 ( );
FILL FILL_32_DFFSR_222 ( );
FILL FILL_33_DFFSR_222 ( );
FILL FILL_34_DFFSR_222 ( );
FILL FILL_35_DFFSR_222 ( );
FILL FILL_36_DFFSR_222 ( );
FILL FILL_37_DFFSR_222 ( );
FILL FILL_38_DFFSR_222 ( );
FILL FILL_39_DFFSR_222 ( );
FILL FILL_40_DFFSR_222 ( );
FILL FILL_41_DFFSR_222 ( );
FILL FILL_42_DFFSR_222 ( );
FILL FILL_43_DFFSR_222 ( );
FILL FILL_44_DFFSR_222 ( );
FILL FILL_45_DFFSR_222 ( );
FILL FILL_46_DFFSR_222 ( );
FILL FILL_47_DFFSR_222 ( );
FILL FILL_48_DFFSR_222 ( );
FILL FILL_49_DFFSR_222 ( );
FILL FILL_50_DFFSR_222 ( );
FILL FILL_0_DFFSR_145 ( );
FILL FILL_1_DFFSR_145 ( );
FILL FILL_2_DFFSR_145 ( );
FILL FILL_3_DFFSR_145 ( );
FILL FILL_4_DFFSR_145 ( );
FILL FILL_5_DFFSR_145 ( );
FILL FILL_6_DFFSR_145 ( );
FILL FILL_7_DFFSR_145 ( );
FILL FILL_8_DFFSR_145 ( );
FILL FILL_9_DFFSR_145 ( );
FILL FILL_10_DFFSR_145 ( );
FILL FILL_11_DFFSR_145 ( );
FILL FILL_12_DFFSR_145 ( );
FILL FILL_13_DFFSR_145 ( );
FILL FILL_14_DFFSR_145 ( );
FILL FILL_15_DFFSR_145 ( );
FILL FILL_16_DFFSR_145 ( );
FILL FILL_17_DFFSR_145 ( );
FILL FILL_18_DFFSR_145 ( );
FILL FILL_19_DFFSR_145 ( );
FILL FILL_20_DFFSR_145 ( );
FILL FILL_21_DFFSR_145 ( );
FILL FILL_22_DFFSR_145 ( );
FILL FILL_23_DFFSR_145 ( );
FILL FILL_24_DFFSR_145 ( );
FILL FILL_25_DFFSR_145 ( );
FILL FILL_26_DFFSR_145 ( );
FILL FILL_27_DFFSR_145 ( );
FILL FILL_28_DFFSR_145 ( );
FILL FILL_29_DFFSR_145 ( );
FILL FILL_30_DFFSR_145 ( );
FILL FILL_31_DFFSR_145 ( );
FILL FILL_32_DFFSR_145 ( );
FILL FILL_33_DFFSR_145 ( );
FILL FILL_34_DFFSR_145 ( );
FILL FILL_35_DFFSR_145 ( );
FILL FILL_36_DFFSR_145 ( );
FILL FILL_37_DFFSR_145 ( );
FILL FILL_38_DFFSR_145 ( );
FILL FILL_39_DFFSR_145 ( );
FILL FILL_40_DFFSR_145 ( );
FILL FILL_41_DFFSR_145 ( );
FILL FILL_42_DFFSR_145 ( );
FILL FILL_43_DFFSR_145 ( );
FILL FILL_44_DFFSR_145 ( );
FILL FILL_45_DFFSR_145 ( );
FILL FILL_46_DFFSR_145 ( );
FILL FILL_47_DFFSR_145 ( );
FILL FILL_48_DFFSR_145 ( );
FILL FILL_49_DFFSR_145 ( );
FILL FILL_50_DFFSR_145 ( );
FILL FILL_0_DFFSR_241 ( );
FILL FILL_1_DFFSR_241 ( );
FILL FILL_2_DFFSR_241 ( );
FILL FILL_3_DFFSR_241 ( );
FILL FILL_4_DFFSR_241 ( );
FILL FILL_5_DFFSR_241 ( );
FILL FILL_6_DFFSR_241 ( );
FILL FILL_7_DFFSR_241 ( );
FILL FILL_8_DFFSR_241 ( );
FILL FILL_9_DFFSR_241 ( );
FILL FILL_10_DFFSR_241 ( );
FILL FILL_11_DFFSR_241 ( );
FILL FILL_12_DFFSR_241 ( );
FILL FILL_13_DFFSR_241 ( );
FILL FILL_14_DFFSR_241 ( );
FILL FILL_15_DFFSR_241 ( );
FILL FILL_16_DFFSR_241 ( );
FILL FILL_17_DFFSR_241 ( );
FILL FILL_18_DFFSR_241 ( );
FILL FILL_19_DFFSR_241 ( );
FILL FILL_20_DFFSR_241 ( );
FILL FILL_21_DFFSR_241 ( );
FILL FILL_22_DFFSR_241 ( );
FILL FILL_23_DFFSR_241 ( );
FILL FILL_24_DFFSR_241 ( );
FILL FILL_25_DFFSR_241 ( );
FILL FILL_26_DFFSR_241 ( );
FILL FILL_27_DFFSR_241 ( );
FILL FILL_28_DFFSR_241 ( );
FILL FILL_29_DFFSR_241 ( );
FILL FILL_30_DFFSR_241 ( );
FILL FILL_31_DFFSR_241 ( );
FILL FILL_32_DFFSR_241 ( );
FILL FILL_33_DFFSR_241 ( );
FILL FILL_34_DFFSR_241 ( );
FILL FILL_35_DFFSR_241 ( );
FILL FILL_36_DFFSR_241 ( );
FILL FILL_37_DFFSR_241 ( );
FILL FILL_38_DFFSR_241 ( );
FILL FILL_39_DFFSR_241 ( );
FILL FILL_40_DFFSR_241 ( );
FILL FILL_41_DFFSR_241 ( );
FILL FILL_42_DFFSR_241 ( );
FILL FILL_43_DFFSR_241 ( );
FILL FILL_44_DFFSR_241 ( );
FILL FILL_45_DFFSR_241 ( );
FILL FILL_46_DFFSR_241 ( );
FILL FILL_47_DFFSR_241 ( );
FILL FILL_48_DFFSR_241 ( );
FILL FILL_49_DFFSR_241 ( );
FILL FILL_50_DFFSR_241 ( );
FILL FILL_0_DFFSR_217 ( );
FILL FILL_1_DFFSR_217 ( );
FILL FILL_2_DFFSR_217 ( );
FILL FILL_3_DFFSR_217 ( );
FILL FILL_4_DFFSR_217 ( );
FILL FILL_5_DFFSR_217 ( );
FILL FILL_6_DFFSR_217 ( );
FILL FILL_7_DFFSR_217 ( );
FILL FILL_8_DFFSR_217 ( );
FILL FILL_9_DFFSR_217 ( );
FILL FILL_10_DFFSR_217 ( );
FILL FILL_11_DFFSR_217 ( );
FILL FILL_12_DFFSR_217 ( );
FILL FILL_13_DFFSR_217 ( );
FILL FILL_14_DFFSR_217 ( );
FILL FILL_15_DFFSR_217 ( );
FILL FILL_16_DFFSR_217 ( );
FILL FILL_17_DFFSR_217 ( );
FILL FILL_18_DFFSR_217 ( );
FILL FILL_19_DFFSR_217 ( );
FILL FILL_20_DFFSR_217 ( );
FILL FILL_21_DFFSR_217 ( );
FILL FILL_22_DFFSR_217 ( );
FILL FILL_23_DFFSR_217 ( );
FILL FILL_24_DFFSR_217 ( );
FILL FILL_25_DFFSR_217 ( );
FILL FILL_26_DFFSR_217 ( );
FILL FILL_27_DFFSR_217 ( );
FILL FILL_28_DFFSR_217 ( );
FILL FILL_29_DFFSR_217 ( );
FILL FILL_30_DFFSR_217 ( );
FILL FILL_31_DFFSR_217 ( );
FILL FILL_32_DFFSR_217 ( );
FILL FILL_33_DFFSR_217 ( );
FILL FILL_34_DFFSR_217 ( );
FILL FILL_35_DFFSR_217 ( );
FILL FILL_36_DFFSR_217 ( );
FILL FILL_37_DFFSR_217 ( );
FILL FILL_38_DFFSR_217 ( );
FILL FILL_39_DFFSR_217 ( );
FILL FILL_40_DFFSR_217 ( );
FILL FILL_41_DFFSR_217 ( );
FILL FILL_42_DFFSR_217 ( );
FILL FILL_43_DFFSR_217 ( );
FILL FILL_44_DFFSR_217 ( );
FILL FILL_45_DFFSR_217 ( );
FILL FILL_46_DFFSR_217 ( );
FILL FILL_47_DFFSR_217 ( );
FILL FILL_48_DFFSR_217 ( );
FILL FILL_49_DFFSR_217 ( );
FILL FILL_50_DFFSR_217 ( );
FILL FILL_51_DFFSR_217 ( );
FILL FILL_0_CLKBUF1_34 ( );
FILL FILL_1_CLKBUF1_34 ( );
FILL FILL_2_CLKBUF1_34 ( );
FILL FILL_3_CLKBUF1_34 ( );
FILL FILL_4_CLKBUF1_34 ( );
FILL FILL_5_CLKBUF1_34 ( );
FILL FILL_6_CLKBUF1_34 ( );
FILL FILL_7_CLKBUF1_34 ( );
FILL FILL_8_CLKBUF1_34 ( );
FILL FILL_9_CLKBUF1_34 ( );
FILL FILL_10_CLKBUF1_34 ( );
FILL FILL_11_CLKBUF1_34 ( );
FILL FILL_12_CLKBUF1_34 ( );
FILL FILL_13_CLKBUF1_34 ( );
FILL FILL_14_CLKBUF1_34 ( );
FILL FILL_15_CLKBUF1_34 ( );
FILL FILL_16_CLKBUF1_34 ( );
FILL FILL_17_CLKBUF1_34 ( );
FILL FILL_18_CLKBUF1_34 ( );
FILL FILL_19_CLKBUF1_34 ( );
FILL FILL_20_CLKBUF1_34 ( );
FILL FILL_0_DFFSR_165 ( );
FILL FILL_1_DFFSR_165 ( );
FILL FILL_2_DFFSR_165 ( );
FILL FILL_3_DFFSR_165 ( );
FILL FILL_4_DFFSR_165 ( );
FILL FILL_5_DFFSR_165 ( );
FILL FILL_6_DFFSR_165 ( );
FILL FILL_7_DFFSR_165 ( );
FILL FILL_8_DFFSR_165 ( );
FILL FILL_9_DFFSR_165 ( );
FILL FILL_10_DFFSR_165 ( );
FILL FILL_11_DFFSR_165 ( );
FILL FILL_12_DFFSR_165 ( );
FILL FILL_13_DFFSR_165 ( );
FILL FILL_14_DFFSR_165 ( );
FILL FILL_15_DFFSR_165 ( );
FILL FILL_16_DFFSR_165 ( );
FILL FILL_17_DFFSR_165 ( );
FILL FILL_18_DFFSR_165 ( );
FILL FILL_19_DFFSR_165 ( );
FILL FILL_20_DFFSR_165 ( );
FILL FILL_21_DFFSR_165 ( );
FILL FILL_22_DFFSR_165 ( );
FILL FILL_23_DFFSR_165 ( );
FILL FILL_24_DFFSR_165 ( );
FILL FILL_25_DFFSR_165 ( );
FILL FILL_26_DFFSR_165 ( );
FILL FILL_27_DFFSR_165 ( );
FILL FILL_28_DFFSR_165 ( );
FILL FILL_29_DFFSR_165 ( );
FILL FILL_30_DFFSR_165 ( );
FILL FILL_31_DFFSR_165 ( );
FILL FILL_32_DFFSR_165 ( );
FILL FILL_33_DFFSR_165 ( );
FILL FILL_34_DFFSR_165 ( );
FILL FILL_35_DFFSR_165 ( );
FILL FILL_36_DFFSR_165 ( );
FILL FILL_37_DFFSR_165 ( );
FILL FILL_38_DFFSR_165 ( );
FILL FILL_39_DFFSR_165 ( );
FILL FILL_40_DFFSR_165 ( );
FILL FILL_41_DFFSR_165 ( );
FILL FILL_42_DFFSR_165 ( );
FILL FILL_43_DFFSR_165 ( );
FILL FILL_44_DFFSR_165 ( );
FILL FILL_45_DFFSR_165 ( );
FILL FILL_46_DFFSR_165 ( );
FILL FILL_47_DFFSR_165 ( );
FILL FILL_48_DFFSR_165 ( );
FILL FILL_49_DFFSR_165 ( );
FILL FILL_50_DFFSR_165 ( );
FILL FILL_0_DFFSR_266 ( );
FILL FILL_1_DFFSR_266 ( );
FILL FILL_2_DFFSR_266 ( );
FILL FILL_3_DFFSR_266 ( );
FILL FILL_4_DFFSR_266 ( );
FILL FILL_5_DFFSR_266 ( );
FILL FILL_6_DFFSR_266 ( );
FILL FILL_7_DFFSR_266 ( );
FILL FILL_8_DFFSR_266 ( );
FILL FILL_9_DFFSR_266 ( );
FILL FILL_10_DFFSR_266 ( );
FILL FILL_11_DFFSR_266 ( );
FILL FILL_12_DFFSR_266 ( );
FILL FILL_13_DFFSR_266 ( );
FILL FILL_14_DFFSR_266 ( );
FILL FILL_15_DFFSR_266 ( );
FILL FILL_16_DFFSR_266 ( );
FILL FILL_17_DFFSR_266 ( );
FILL FILL_18_DFFSR_266 ( );
FILL FILL_19_DFFSR_266 ( );
FILL FILL_20_DFFSR_266 ( );
FILL FILL_21_DFFSR_266 ( );
FILL FILL_22_DFFSR_266 ( );
FILL FILL_23_DFFSR_266 ( );
FILL FILL_24_DFFSR_266 ( );
FILL FILL_25_DFFSR_266 ( );
FILL FILL_26_DFFSR_266 ( );
FILL FILL_27_DFFSR_266 ( );
FILL FILL_28_DFFSR_266 ( );
FILL FILL_29_DFFSR_266 ( );
FILL FILL_30_DFFSR_266 ( );
FILL FILL_31_DFFSR_266 ( );
FILL FILL_32_DFFSR_266 ( );
FILL FILL_33_DFFSR_266 ( );
FILL FILL_34_DFFSR_266 ( );
FILL FILL_35_DFFSR_266 ( );
FILL FILL_36_DFFSR_266 ( );
FILL FILL_37_DFFSR_266 ( );
FILL FILL_38_DFFSR_266 ( );
FILL FILL_39_DFFSR_266 ( );
FILL FILL_40_DFFSR_266 ( );
FILL FILL_41_DFFSR_266 ( );
FILL FILL_42_DFFSR_266 ( );
FILL FILL_43_DFFSR_266 ( );
FILL FILL_44_DFFSR_266 ( );
FILL FILL_45_DFFSR_266 ( );
FILL FILL_46_DFFSR_266 ( );
FILL FILL_47_DFFSR_266 ( );
FILL FILL_48_DFFSR_266 ( );
FILL FILL_49_DFFSR_266 ( );
FILL FILL_50_DFFSR_266 ( );
FILL FILL_0_NAND3X1_138 ( );
FILL FILL_1_NAND3X1_138 ( );
FILL FILL_2_NAND3X1_138 ( );
FILL FILL_3_NAND3X1_138 ( );
FILL FILL_4_NAND3X1_138 ( );
FILL FILL_5_NAND3X1_138 ( );
FILL FILL_6_NAND3X1_138 ( );
FILL FILL_7_NAND3X1_138 ( );
FILL FILL_8_NAND3X1_138 ( );
FILL FILL_0_OAI21X1_23 ( );
FILL FILL_1_OAI21X1_23 ( );
FILL FILL_2_OAI21X1_23 ( );
FILL FILL_3_OAI21X1_23 ( );
FILL FILL_4_OAI21X1_23 ( );
FILL FILL_5_OAI21X1_23 ( );
FILL FILL_6_OAI21X1_23 ( );
FILL FILL_7_OAI21X1_23 ( );
FILL FILL_8_OAI21X1_23 ( );
FILL FILL_0_INVX1_141 ( );
FILL FILL_1_INVX1_141 ( );
FILL FILL_2_INVX1_141 ( );
FILL FILL_3_INVX1_141 ( );
FILL FILL_0_DFFSR_269 ( );
FILL FILL_1_DFFSR_269 ( );
FILL FILL_2_DFFSR_269 ( );
FILL FILL_3_DFFSR_269 ( );
FILL FILL_4_DFFSR_269 ( );
FILL FILL_5_DFFSR_269 ( );
FILL FILL_6_DFFSR_269 ( );
FILL FILL_7_DFFSR_269 ( );
FILL FILL_8_DFFSR_269 ( );
FILL FILL_9_DFFSR_269 ( );
FILL FILL_10_DFFSR_269 ( );
FILL FILL_11_DFFSR_269 ( );
FILL FILL_12_DFFSR_269 ( );
FILL FILL_13_DFFSR_269 ( );
FILL FILL_14_DFFSR_269 ( );
FILL FILL_15_DFFSR_269 ( );
FILL FILL_16_DFFSR_269 ( );
FILL FILL_17_DFFSR_269 ( );
FILL FILL_18_DFFSR_269 ( );
FILL FILL_19_DFFSR_269 ( );
FILL FILL_20_DFFSR_269 ( );
FILL FILL_21_DFFSR_269 ( );
FILL FILL_22_DFFSR_269 ( );
FILL FILL_23_DFFSR_269 ( );
FILL FILL_24_DFFSR_269 ( );
FILL FILL_25_DFFSR_269 ( );
FILL FILL_26_DFFSR_269 ( );
FILL FILL_27_DFFSR_269 ( );
FILL FILL_28_DFFSR_269 ( );
FILL FILL_29_DFFSR_269 ( );
FILL FILL_30_DFFSR_269 ( );
FILL FILL_31_DFFSR_269 ( );
FILL FILL_32_DFFSR_269 ( );
FILL FILL_33_DFFSR_269 ( );
FILL FILL_34_DFFSR_269 ( );
FILL FILL_35_DFFSR_269 ( );
FILL FILL_36_DFFSR_269 ( );
FILL FILL_37_DFFSR_269 ( );
FILL FILL_38_DFFSR_269 ( );
FILL FILL_39_DFFSR_269 ( );
FILL FILL_40_DFFSR_269 ( );
FILL FILL_41_DFFSR_269 ( );
FILL FILL_42_DFFSR_269 ( );
FILL FILL_43_DFFSR_269 ( );
FILL FILL_44_DFFSR_269 ( );
FILL FILL_45_DFFSR_269 ( );
FILL FILL_46_DFFSR_269 ( );
FILL FILL_47_DFFSR_269 ( );
FILL FILL_48_DFFSR_269 ( );
FILL FILL_49_DFFSR_269 ( );
FILL FILL_50_DFFSR_269 ( );
FILL FILL_0_AOI21X1_57 ( );
FILL FILL_1_AOI21X1_57 ( );
FILL FILL_2_AOI21X1_57 ( );
FILL FILL_3_AOI21X1_57 ( );
FILL FILL_4_AOI21X1_57 ( );
FILL FILL_5_AOI21X1_57 ( );
FILL FILL_6_AOI21X1_57 ( );
FILL FILL_7_AOI21X1_57 ( );
FILL FILL_8_AOI21X1_57 ( );
FILL FILL_0_NAND2X1_163 ( );
FILL FILL_1_NAND2X1_163 ( );
FILL FILL_2_NAND2X1_163 ( );
FILL FILL_3_NAND2X1_163 ( );
FILL FILL_4_NAND2X1_163 ( );
FILL FILL_5_NAND2X1_163 ( );
FILL FILL_6_NAND2X1_163 ( );
FILL FILL_0_NAND2X1_143 ( );
FILL FILL_1_NAND2X1_143 ( );
FILL FILL_2_NAND2X1_143 ( );
FILL FILL_3_NAND2X1_143 ( );
FILL FILL_4_NAND2X1_143 ( );
FILL FILL_5_NAND2X1_143 ( );
FILL FILL_6_NAND2X1_143 ( );
FILL FILL_0_OAI21X1_104 ( );
FILL FILL_1_OAI21X1_104 ( );
FILL FILL_2_OAI21X1_104 ( );
FILL FILL_3_OAI21X1_104 ( );
FILL FILL_4_OAI21X1_104 ( );
FILL FILL_5_OAI21X1_104 ( );
FILL FILL_6_OAI21X1_104 ( );
FILL FILL_7_OAI21X1_104 ( );
FILL FILL_8_OAI21X1_104 ( );
FILL FILL_0_DFFPOSX1_32 ( );
FILL FILL_1_DFFPOSX1_32 ( );
FILL FILL_2_DFFPOSX1_32 ( );
FILL FILL_3_DFFPOSX1_32 ( );
FILL FILL_4_DFFPOSX1_32 ( );
FILL FILL_5_DFFPOSX1_32 ( );
FILL FILL_6_DFFPOSX1_32 ( );
FILL FILL_7_DFFPOSX1_32 ( );
FILL FILL_8_DFFPOSX1_32 ( );
FILL FILL_9_DFFPOSX1_32 ( );
FILL FILL_10_DFFPOSX1_32 ( );
FILL FILL_11_DFFPOSX1_32 ( );
FILL FILL_12_DFFPOSX1_32 ( );
FILL FILL_13_DFFPOSX1_32 ( );
FILL FILL_14_DFFPOSX1_32 ( );
FILL FILL_15_DFFPOSX1_32 ( );
FILL FILL_16_DFFPOSX1_32 ( );
FILL FILL_17_DFFPOSX1_32 ( );
FILL FILL_18_DFFPOSX1_32 ( );
FILL FILL_19_DFFPOSX1_32 ( );
FILL FILL_20_DFFPOSX1_32 ( );
FILL FILL_21_DFFPOSX1_32 ( );
FILL FILL_22_DFFPOSX1_32 ( );
FILL FILL_23_DFFPOSX1_32 ( );
FILL FILL_24_DFFPOSX1_32 ( );
FILL FILL_25_DFFPOSX1_32 ( );
FILL FILL_26_DFFPOSX1_32 ( );
FILL FILL_27_DFFPOSX1_32 ( );
FILL FILL_0_NOR2X1_62 ( );
FILL FILL_1_NOR2X1_62 ( );
FILL FILL_2_NOR2X1_62 ( );
FILL FILL_3_NOR2X1_62 ( );
FILL FILL_4_NOR2X1_62 ( );
FILL FILL_5_NOR2X1_62 ( );
FILL FILL_6_NOR2X1_62 ( );
FILL FILL_0_DFFPOSX1_10 ( );
FILL FILL_1_DFFPOSX1_10 ( );
FILL FILL_2_DFFPOSX1_10 ( );
FILL FILL_3_DFFPOSX1_10 ( );
FILL FILL_4_DFFPOSX1_10 ( );
FILL FILL_5_DFFPOSX1_10 ( );
FILL FILL_6_DFFPOSX1_10 ( );
FILL FILL_7_DFFPOSX1_10 ( );
FILL FILL_8_DFFPOSX1_10 ( );
FILL FILL_9_DFFPOSX1_10 ( );
FILL FILL_10_DFFPOSX1_10 ( );
FILL FILL_11_DFFPOSX1_10 ( );
FILL FILL_12_DFFPOSX1_10 ( );
FILL FILL_13_DFFPOSX1_10 ( );
FILL FILL_14_DFFPOSX1_10 ( );
FILL FILL_15_DFFPOSX1_10 ( );
FILL FILL_16_DFFPOSX1_10 ( );
FILL FILL_17_DFFPOSX1_10 ( );
FILL FILL_18_DFFPOSX1_10 ( );
FILL FILL_19_DFFPOSX1_10 ( );
FILL FILL_20_DFFPOSX1_10 ( );
FILL FILL_21_DFFPOSX1_10 ( );
FILL FILL_22_DFFPOSX1_10 ( );
FILL FILL_23_DFFPOSX1_10 ( );
FILL FILL_24_DFFPOSX1_10 ( );
FILL FILL_25_DFFPOSX1_10 ( );
FILL FILL_26_DFFPOSX1_10 ( );
FILL FILL_27_DFFPOSX1_10 ( );
FILL FILL_0_CLKBUF1_25 ( );
FILL FILL_1_CLKBUF1_25 ( );
FILL FILL_2_CLKBUF1_25 ( );
FILL FILL_3_CLKBUF1_25 ( );
FILL FILL_4_CLKBUF1_25 ( );
FILL FILL_5_CLKBUF1_25 ( );
FILL FILL_6_CLKBUF1_25 ( );
FILL FILL_7_CLKBUF1_25 ( );
FILL FILL_8_CLKBUF1_25 ( );
FILL FILL_9_CLKBUF1_25 ( );
FILL FILL_10_CLKBUF1_25 ( );
FILL FILL_11_CLKBUF1_25 ( );
FILL FILL_12_CLKBUF1_25 ( );
FILL FILL_13_CLKBUF1_25 ( );
FILL FILL_14_CLKBUF1_25 ( );
FILL FILL_15_CLKBUF1_25 ( );
FILL FILL_16_CLKBUF1_25 ( );
FILL FILL_17_CLKBUF1_25 ( );
FILL FILL_18_CLKBUF1_25 ( );
FILL FILL_19_CLKBUF1_25 ( );
FILL FILL_20_CLKBUF1_25 ( );
FILL FILL_0_DFFSR_230 ( );
FILL FILL_1_DFFSR_230 ( );
FILL FILL_2_DFFSR_230 ( );
FILL FILL_3_DFFSR_230 ( );
FILL FILL_4_DFFSR_230 ( );
FILL FILL_5_DFFSR_230 ( );
FILL FILL_6_DFFSR_230 ( );
FILL FILL_7_DFFSR_230 ( );
FILL FILL_8_DFFSR_230 ( );
FILL FILL_9_DFFSR_230 ( );
FILL FILL_10_DFFSR_230 ( );
FILL FILL_11_DFFSR_230 ( );
FILL FILL_12_DFFSR_230 ( );
FILL FILL_13_DFFSR_230 ( );
FILL FILL_14_DFFSR_230 ( );
FILL FILL_15_DFFSR_230 ( );
FILL FILL_16_DFFSR_230 ( );
FILL FILL_17_DFFSR_230 ( );
FILL FILL_18_DFFSR_230 ( );
FILL FILL_19_DFFSR_230 ( );
FILL FILL_20_DFFSR_230 ( );
FILL FILL_21_DFFSR_230 ( );
FILL FILL_22_DFFSR_230 ( );
FILL FILL_23_DFFSR_230 ( );
FILL FILL_24_DFFSR_230 ( );
FILL FILL_25_DFFSR_230 ( );
FILL FILL_26_DFFSR_230 ( );
FILL FILL_27_DFFSR_230 ( );
FILL FILL_28_DFFSR_230 ( );
FILL FILL_29_DFFSR_230 ( );
FILL FILL_30_DFFSR_230 ( );
FILL FILL_31_DFFSR_230 ( );
FILL FILL_32_DFFSR_230 ( );
FILL FILL_33_DFFSR_230 ( );
FILL FILL_34_DFFSR_230 ( );
FILL FILL_35_DFFSR_230 ( );
FILL FILL_36_DFFSR_230 ( );
FILL FILL_37_DFFSR_230 ( );
FILL FILL_38_DFFSR_230 ( );
FILL FILL_39_DFFSR_230 ( );
FILL FILL_40_DFFSR_230 ( );
FILL FILL_41_DFFSR_230 ( );
FILL FILL_42_DFFSR_230 ( );
FILL FILL_43_DFFSR_230 ( );
FILL FILL_44_DFFSR_230 ( );
FILL FILL_45_DFFSR_230 ( );
FILL FILL_46_DFFSR_230 ( );
FILL FILL_47_DFFSR_230 ( );
FILL FILL_48_DFFSR_230 ( );
FILL FILL_49_DFFSR_230 ( );
FILL FILL_50_DFFSR_230 ( );
FILL FILL_0_DFFPOSX1_9 ( );
FILL FILL_1_DFFPOSX1_9 ( );
FILL FILL_2_DFFPOSX1_9 ( );
FILL FILL_3_DFFPOSX1_9 ( );
FILL FILL_4_DFFPOSX1_9 ( );
FILL FILL_5_DFFPOSX1_9 ( );
FILL FILL_6_DFFPOSX1_9 ( );
FILL FILL_7_DFFPOSX1_9 ( );
FILL FILL_8_DFFPOSX1_9 ( );
FILL FILL_9_DFFPOSX1_9 ( );
FILL FILL_10_DFFPOSX1_9 ( );
FILL FILL_11_DFFPOSX1_9 ( );
FILL FILL_12_DFFPOSX1_9 ( );
FILL FILL_13_DFFPOSX1_9 ( );
FILL FILL_14_DFFPOSX1_9 ( );
FILL FILL_15_DFFPOSX1_9 ( );
FILL FILL_16_DFFPOSX1_9 ( );
FILL FILL_17_DFFPOSX1_9 ( );
FILL FILL_18_DFFPOSX1_9 ( );
FILL FILL_19_DFFPOSX1_9 ( );
FILL FILL_20_DFFPOSX1_9 ( );
FILL FILL_21_DFFPOSX1_9 ( );
FILL FILL_22_DFFPOSX1_9 ( );
FILL FILL_23_DFFPOSX1_9 ( );
FILL FILL_24_DFFPOSX1_9 ( );
FILL FILL_25_DFFPOSX1_9 ( );
FILL FILL_26_DFFPOSX1_9 ( );
FILL FILL_27_DFFPOSX1_9 ( );
FILL FILL_0_DFFSR_153 ( );
FILL FILL_1_DFFSR_153 ( );
FILL FILL_2_DFFSR_153 ( );
FILL FILL_3_DFFSR_153 ( );
FILL FILL_4_DFFSR_153 ( );
FILL FILL_5_DFFSR_153 ( );
FILL FILL_6_DFFSR_153 ( );
FILL FILL_7_DFFSR_153 ( );
FILL FILL_8_DFFSR_153 ( );
FILL FILL_9_DFFSR_153 ( );
FILL FILL_10_DFFSR_153 ( );
FILL FILL_11_DFFSR_153 ( );
FILL FILL_12_DFFSR_153 ( );
FILL FILL_13_DFFSR_153 ( );
FILL FILL_14_DFFSR_153 ( );
FILL FILL_15_DFFSR_153 ( );
FILL FILL_16_DFFSR_153 ( );
FILL FILL_17_DFFSR_153 ( );
FILL FILL_18_DFFSR_153 ( );
FILL FILL_19_DFFSR_153 ( );
FILL FILL_20_DFFSR_153 ( );
FILL FILL_21_DFFSR_153 ( );
FILL FILL_22_DFFSR_153 ( );
FILL FILL_23_DFFSR_153 ( );
FILL FILL_24_DFFSR_153 ( );
FILL FILL_25_DFFSR_153 ( );
FILL FILL_26_DFFSR_153 ( );
FILL FILL_27_DFFSR_153 ( );
FILL FILL_28_DFFSR_153 ( );
FILL FILL_29_DFFSR_153 ( );
FILL FILL_30_DFFSR_153 ( );
FILL FILL_31_DFFSR_153 ( );
FILL FILL_32_DFFSR_153 ( );
FILL FILL_33_DFFSR_153 ( );
FILL FILL_34_DFFSR_153 ( );
FILL FILL_35_DFFSR_153 ( );
FILL FILL_36_DFFSR_153 ( );
FILL FILL_37_DFFSR_153 ( );
FILL FILL_38_DFFSR_153 ( );
FILL FILL_39_DFFSR_153 ( );
FILL FILL_40_DFFSR_153 ( );
FILL FILL_41_DFFSR_153 ( );
FILL FILL_42_DFFSR_153 ( );
FILL FILL_43_DFFSR_153 ( );
FILL FILL_44_DFFSR_153 ( );
FILL FILL_45_DFFSR_153 ( );
FILL FILL_46_DFFSR_153 ( );
FILL FILL_47_DFFSR_153 ( );
FILL FILL_48_DFFSR_153 ( );
FILL FILL_49_DFFSR_153 ( );
FILL FILL_50_DFFSR_153 ( );
FILL FILL_0_INVX1_67 ( );
FILL FILL_1_INVX1_67 ( );
FILL FILL_2_INVX1_67 ( );
FILL FILL_3_INVX1_67 ( );
FILL FILL_4_INVX1_67 ( );
FILL FILL_0_NAND2X1_35 ( );
FILL FILL_1_NAND2X1_35 ( );
FILL FILL_2_NAND2X1_35 ( );
FILL FILL_3_NAND2X1_35 ( );
FILL FILL_4_NAND2X1_35 ( );
FILL FILL_5_NAND2X1_35 ( );
FILL FILL_6_NAND2X1_35 ( );
FILL FILL_0_INVX1_68 ( );
FILL FILL_1_INVX1_68 ( );
FILL FILL_2_INVX1_68 ( );
FILL FILL_3_INVX1_68 ( );
FILL FILL_4_INVX1_68 ( );
FILL FILL_0_OAI21X1_9 ( );
FILL FILL_1_OAI21X1_9 ( );
FILL FILL_2_OAI21X1_9 ( );
FILL FILL_3_OAI21X1_9 ( );
FILL FILL_4_OAI21X1_9 ( );
FILL FILL_5_OAI21X1_9 ( );
FILL FILL_6_OAI21X1_9 ( );
FILL FILL_7_OAI21X1_9 ( );
FILL FILL_8_OAI21X1_9 ( );
FILL FILL_9_OAI21X1_9 ( );
FILL FILL_0_INVX1_106 ( );
FILL FILL_1_INVX1_106 ( );
FILL FILL_2_INVX1_106 ( );
FILL FILL_3_INVX1_106 ( );
FILL FILL_0_DFFSR_201 ( );
FILL FILL_1_DFFSR_201 ( );
FILL FILL_2_DFFSR_201 ( );
FILL FILL_3_DFFSR_201 ( );
FILL FILL_4_DFFSR_201 ( );
FILL FILL_5_DFFSR_201 ( );
FILL FILL_6_DFFSR_201 ( );
FILL FILL_7_DFFSR_201 ( );
FILL FILL_8_DFFSR_201 ( );
FILL FILL_9_DFFSR_201 ( );
FILL FILL_10_DFFSR_201 ( );
FILL FILL_11_DFFSR_201 ( );
FILL FILL_12_DFFSR_201 ( );
FILL FILL_13_DFFSR_201 ( );
FILL FILL_14_DFFSR_201 ( );
FILL FILL_15_DFFSR_201 ( );
FILL FILL_16_DFFSR_201 ( );
FILL FILL_17_DFFSR_201 ( );
FILL FILL_18_DFFSR_201 ( );
FILL FILL_19_DFFSR_201 ( );
FILL FILL_20_DFFSR_201 ( );
FILL FILL_21_DFFSR_201 ( );
FILL FILL_22_DFFSR_201 ( );
FILL FILL_23_DFFSR_201 ( );
FILL FILL_24_DFFSR_201 ( );
FILL FILL_25_DFFSR_201 ( );
FILL FILL_26_DFFSR_201 ( );
FILL FILL_27_DFFSR_201 ( );
FILL FILL_28_DFFSR_201 ( );
FILL FILL_29_DFFSR_201 ( );
FILL FILL_30_DFFSR_201 ( );
FILL FILL_31_DFFSR_201 ( );
FILL FILL_32_DFFSR_201 ( );
FILL FILL_33_DFFSR_201 ( );
FILL FILL_34_DFFSR_201 ( );
FILL FILL_35_DFFSR_201 ( );
FILL FILL_36_DFFSR_201 ( );
FILL FILL_37_DFFSR_201 ( );
FILL FILL_38_DFFSR_201 ( );
FILL FILL_39_DFFSR_201 ( );
FILL FILL_40_DFFSR_201 ( );
FILL FILL_41_DFFSR_201 ( );
FILL FILL_42_DFFSR_201 ( );
FILL FILL_43_DFFSR_201 ( );
FILL FILL_44_DFFSR_201 ( );
FILL FILL_45_DFFSR_201 ( );
FILL FILL_46_DFFSR_201 ( );
FILL FILL_47_DFFSR_201 ( );
FILL FILL_48_DFFSR_201 ( );
FILL FILL_49_DFFSR_201 ( );
FILL FILL_50_DFFSR_201 ( );
FILL FILL_0_INVX1_94 ( );
FILL FILL_1_INVX1_94 ( );
FILL FILL_2_INVX1_94 ( );
FILL FILL_3_INVX1_94 ( );
FILL FILL_4_INVX1_94 ( );
FILL FILL_0_CLKBUF1_10 ( );
FILL FILL_1_CLKBUF1_10 ( );
FILL FILL_2_CLKBUF1_10 ( );
FILL FILL_3_CLKBUF1_10 ( );
FILL FILL_4_CLKBUF1_10 ( );
FILL FILL_5_CLKBUF1_10 ( );
FILL FILL_6_CLKBUF1_10 ( );
FILL FILL_7_CLKBUF1_10 ( );
FILL FILL_8_CLKBUF1_10 ( );
FILL FILL_9_CLKBUF1_10 ( );
FILL FILL_10_CLKBUF1_10 ( );
FILL FILL_11_CLKBUF1_10 ( );
FILL FILL_12_CLKBUF1_10 ( );
FILL FILL_13_CLKBUF1_10 ( );
FILL FILL_14_CLKBUF1_10 ( );
FILL FILL_15_CLKBUF1_10 ( );
FILL FILL_16_CLKBUF1_10 ( );
FILL FILL_17_CLKBUF1_10 ( );
FILL FILL_18_CLKBUF1_10 ( );
FILL FILL_19_CLKBUF1_10 ( );
FILL FILL_0_OAI21X1_94 ( );
FILL FILL_1_OAI21X1_94 ( );
FILL FILL_2_OAI21X1_94 ( );
FILL FILL_3_OAI21X1_94 ( );
FILL FILL_4_OAI21X1_94 ( );
FILL FILL_5_OAI21X1_94 ( );
FILL FILL_6_OAI21X1_94 ( );
FILL FILL_7_OAI21X1_94 ( );
FILL FILL_8_OAI21X1_94 ( );
FILL FILL_9_OAI21X1_94 ( );
FILL FILL_0_INVX1_191 ( );
FILL FILL_1_INVX1_191 ( );
FILL FILL_2_INVX1_191 ( );
FILL FILL_3_INVX1_191 ( );
FILL FILL_0_DFFSR_265 ( );
FILL FILL_1_DFFSR_265 ( );
FILL FILL_2_DFFSR_265 ( );
FILL FILL_3_DFFSR_265 ( );
FILL FILL_4_DFFSR_265 ( );
FILL FILL_5_DFFSR_265 ( );
FILL FILL_6_DFFSR_265 ( );
FILL FILL_7_DFFSR_265 ( );
FILL FILL_8_DFFSR_265 ( );
FILL FILL_9_DFFSR_265 ( );
FILL FILL_10_DFFSR_265 ( );
FILL FILL_11_DFFSR_265 ( );
FILL FILL_12_DFFSR_265 ( );
FILL FILL_13_DFFSR_265 ( );
FILL FILL_14_DFFSR_265 ( );
FILL FILL_15_DFFSR_265 ( );
FILL FILL_16_DFFSR_265 ( );
FILL FILL_17_DFFSR_265 ( );
FILL FILL_18_DFFSR_265 ( );
FILL FILL_19_DFFSR_265 ( );
FILL FILL_20_DFFSR_265 ( );
FILL FILL_21_DFFSR_265 ( );
FILL FILL_22_DFFSR_265 ( );
FILL FILL_23_DFFSR_265 ( );
FILL FILL_24_DFFSR_265 ( );
FILL FILL_25_DFFSR_265 ( );
FILL FILL_26_DFFSR_265 ( );
FILL FILL_27_DFFSR_265 ( );
FILL FILL_28_DFFSR_265 ( );
FILL FILL_29_DFFSR_265 ( );
FILL FILL_30_DFFSR_265 ( );
FILL FILL_31_DFFSR_265 ( );
FILL FILL_32_DFFSR_265 ( );
FILL FILL_33_DFFSR_265 ( );
FILL FILL_34_DFFSR_265 ( );
FILL FILL_35_DFFSR_265 ( );
FILL FILL_36_DFFSR_265 ( );
FILL FILL_37_DFFSR_265 ( );
FILL FILL_38_DFFSR_265 ( );
FILL FILL_39_DFFSR_265 ( );
FILL FILL_40_DFFSR_265 ( );
FILL FILL_41_DFFSR_265 ( );
FILL FILL_42_DFFSR_265 ( );
FILL FILL_43_DFFSR_265 ( );
FILL FILL_44_DFFSR_265 ( );
FILL FILL_45_DFFSR_265 ( );
FILL FILL_46_DFFSR_265 ( );
FILL FILL_47_DFFSR_265 ( );
FILL FILL_48_DFFSR_265 ( );
FILL FILL_49_DFFSR_265 ( );
FILL FILL_50_DFFSR_265 ( );
FILL FILL_51_DFFSR_265 ( );
FILL FILL_0_AOI21X1_16 ( );
FILL FILL_1_AOI21X1_16 ( );
FILL FILL_2_AOI21X1_16 ( );
FILL FILL_3_AOI21X1_16 ( );
FILL FILL_4_AOI21X1_16 ( );
FILL FILL_5_AOI21X1_16 ( );
FILL FILL_6_AOI21X1_16 ( );
FILL FILL_7_AOI21X1_16 ( );
FILL FILL_8_AOI21X1_16 ( );
FILL FILL_0_INVX1_153 ( );
FILL FILL_1_INVX1_153 ( );
FILL FILL_2_INVX1_153 ( );
FILL FILL_3_INVX1_153 ( );
FILL FILL_4_INVX1_153 ( );
FILL FILL_0_NOR2X1_67 ( );
FILL FILL_1_NOR2X1_67 ( );
FILL FILL_2_NOR2X1_67 ( );
FILL FILL_3_NOR2X1_67 ( );
FILL FILL_4_NOR2X1_67 ( );
FILL FILL_5_NOR2X1_67 ( );
FILL FILL_6_NOR2X1_67 ( );
FILL FILL_0_NAND3X1_142 ( );
FILL FILL_1_NAND3X1_142 ( );
FILL FILL_2_NAND3X1_142 ( );
FILL FILL_3_NAND3X1_142 ( );
FILL FILL_4_NAND3X1_142 ( );
FILL FILL_5_NAND3X1_142 ( );
FILL FILL_6_NAND3X1_142 ( );
FILL FILL_7_NAND3X1_142 ( );
FILL FILL_8_NAND3X1_142 ( );
FILL FILL_9_NAND3X1_142 ( );
FILL FILL_0_DFFPOSX1_16 ( );
FILL FILL_1_DFFPOSX1_16 ( );
FILL FILL_2_DFFPOSX1_16 ( );
FILL FILL_3_DFFPOSX1_16 ( );
FILL FILL_4_DFFPOSX1_16 ( );
FILL FILL_5_DFFPOSX1_16 ( );
FILL FILL_6_DFFPOSX1_16 ( );
FILL FILL_7_DFFPOSX1_16 ( );
FILL FILL_8_DFFPOSX1_16 ( );
FILL FILL_9_DFFPOSX1_16 ( );
FILL FILL_10_DFFPOSX1_16 ( );
FILL FILL_11_DFFPOSX1_16 ( );
FILL FILL_12_DFFPOSX1_16 ( );
FILL FILL_13_DFFPOSX1_16 ( );
FILL FILL_14_DFFPOSX1_16 ( );
FILL FILL_15_DFFPOSX1_16 ( );
FILL FILL_16_DFFPOSX1_16 ( );
FILL FILL_17_DFFPOSX1_16 ( );
FILL FILL_18_DFFPOSX1_16 ( );
FILL FILL_19_DFFPOSX1_16 ( );
FILL FILL_20_DFFPOSX1_16 ( );
FILL FILL_21_DFFPOSX1_16 ( );
FILL FILL_22_DFFPOSX1_16 ( );
FILL FILL_23_DFFPOSX1_16 ( );
FILL FILL_24_DFFPOSX1_16 ( );
FILL FILL_25_DFFPOSX1_16 ( );
FILL FILL_26_DFFPOSX1_16 ( );
FILL FILL_27_DFFPOSX1_16 ( );
FILL FILL_0_NAND2X1_164 ( );
FILL FILL_1_NAND2X1_164 ( );
FILL FILL_2_NAND2X1_164 ( );
FILL FILL_3_NAND2X1_164 ( );
FILL FILL_4_NAND2X1_164 ( );
FILL FILL_5_NAND2X1_164 ( );
FILL FILL_6_NAND2X1_164 ( );
FILL FILL_0_NAND2X1_142 ( );
FILL FILL_1_NAND2X1_142 ( );
FILL FILL_2_NAND2X1_142 ( );
FILL FILL_3_NAND2X1_142 ( );
FILL FILL_4_NAND2X1_142 ( );
FILL FILL_5_NAND2X1_142 ( );
FILL FILL_6_NAND2X1_142 ( );
FILL FILL_0_AOI21X1_47 ( );
FILL FILL_1_AOI21X1_47 ( );
FILL FILL_2_AOI21X1_47 ( );
FILL FILL_3_AOI21X1_47 ( );
FILL FILL_4_AOI21X1_47 ( );
FILL FILL_5_AOI21X1_47 ( );
FILL FILL_6_AOI21X1_47 ( );
FILL FILL_7_AOI21X1_47 ( );
FILL FILL_8_AOI21X1_47 ( );
FILL FILL_9_AOI21X1_47 ( );
FILL FILL_0_NAND2X1_148 ( );
FILL FILL_1_NAND2X1_148 ( );
FILL FILL_2_NAND2X1_148 ( );
FILL FILL_3_NAND2X1_148 ( );
FILL FILL_4_NAND2X1_148 ( );
FILL FILL_5_NAND2X1_148 ( );
FILL FILL_6_NAND2X1_148 ( );
FILL FILL_0_AOI21X1_50 ( );
FILL FILL_1_AOI21X1_50 ( );
FILL FILL_2_AOI21X1_50 ( );
FILL FILL_3_AOI21X1_50 ( );
FILL FILL_4_AOI21X1_50 ( );
FILL FILL_5_AOI21X1_50 ( );
FILL FILL_6_AOI21X1_50 ( );
FILL FILL_7_AOI21X1_50 ( );
FILL FILL_8_AOI21X1_50 ( );
FILL FILL_9_AOI21X1_50 ( );
FILL FILL_0_NAND2X1_122 ( );
FILL FILL_1_NAND2X1_122 ( );
FILL FILL_2_NAND2X1_122 ( );
FILL FILL_3_NAND2X1_122 ( );
FILL FILL_4_NAND2X1_122 ( );
FILL FILL_5_NAND2X1_122 ( );
FILL FILL_6_NAND2X1_122 ( );
FILL FILL_0_DFFSR_148 ( );
FILL FILL_1_DFFSR_148 ( );
FILL FILL_2_DFFSR_148 ( );
FILL FILL_3_DFFSR_148 ( );
FILL FILL_4_DFFSR_148 ( );
FILL FILL_5_DFFSR_148 ( );
FILL FILL_6_DFFSR_148 ( );
FILL FILL_7_DFFSR_148 ( );
FILL FILL_8_DFFSR_148 ( );
FILL FILL_9_DFFSR_148 ( );
FILL FILL_10_DFFSR_148 ( );
FILL FILL_11_DFFSR_148 ( );
FILL FILL_12_DFFSR_148 ( );
FILL FILL_13_DFFSR_148 ( );
FILL FILL_14_DFFSR_148 ( );
FILL FILL_15_DFFSR_148 ( );
FILL FILL_16_DFFSR_148 ( );
FILL FILL_17_DFFSR_148 ( );
FILL FILL_18_DFFSR_148 ( );
FILL FILL_19_DFFSR_148 ( );
FILL FILL_20_DFFSR_148 ( );
FILL FILL_21_DFFSR_148 ( );
FILL FILL_22_DFFSR_148 ( );
FILL FILL_23_DFFSR_148 ( );
FILL FILL_24_DFFSR_148 ( );
FILL FILL_25_DFFSR_148 ( );
FILL FILL_26_DFFSR_148 ( );
FILL FILL_27_DFFSR_148 ( );
FILL FILL_28_DFFSR_148 ( );
FILL FILL_29_DFFSR_148 ( );
FILL FILL_30_DFFSR_148 ( );
FILL FILL_31_DFFSR_148 ( );
FILL FILL_32_DFFSR_148 ( );
FILL FILL_33_DFFSR_148 ( );
FILL FILL_34_DFFSR_148 ( );
FILL FILL_35_DFFSR_148 ( );
FILL FILL_36_DFFSR_148 ( );
FILL FILL_37_DFFSR_148 ( );
FILL FILL_38_DFFSR_148 ( );
FILL FILL_39_DFFSR_148 ( );
FILL FILL_40_DFFSR_148 ( );
FILL FILL_41_DFFSR_148 ( );
FILL FILL_42_DFFSR_148 ( );
FILL FILL_43_DFFSR_148 ( );
FILL FILL_44_DFFSR_148 ( );
FILL FILL_45_DFFSR_148 ( );
FILL FILL_46_DFFSR_148 ( );
FILL FILL_47_DFFSR_148 ( );
FILL FILL_48_DFFSR_148 ( );
FILL FILL_49_DFFSR_148 ( );
FILL FILL_50_DFFSR_148 ( );
FILL FILL_0_DFFSR_219 ( );
FILL FILL_1_DFFSR_219 ( );
FILL FILL_2_DFFSR_219 ( );
FILL FILL_3_DFFSR_219 ( );
FILL FILL_4_DFFSR_219 ( );
FILL FILL_5_DFFSR_219 ( );
FILL FILL_6_DFFSR_219 ( );
FILL FILL_7_DFFSR_219 ( );
FILL FILL_8_DFFSR_219 ( );
FILL FILL_9_DFFSR_219 ( );
FILL FILL_10_DFFSR_219 ( );
FILL FILL_11_DFFSR_219 ( );
FILL FILL_12_DFFSR_219 ( );
FILL FILL_13_DFFSR_219 ( );
FILL FILL_14_DFFSR_219 ( );
FILL FILL_15_DFFSR_219 ( );
FILL FILL_16_DFFSR_219 ( );
FILL FILL_17_DFFSR_219 ( );
FILL FILL_18_DFFSR_219 ( );
FILL FILL_19_DFFSR_219 ( );
FILL FILL_20_DFFSR_219 ( );
FILL FILL_21_DFFSR_219 ( );
FILL FILL_22_DFFSR_219 ( );
FILL FILL_23_DFFSR_219 ( );
FILL FILL_24_DFFSR_219 ( );
FILL FILL_25_DFFSR_219 ( );
FILL FILL_26_DFFSR_219 ( );
FILL FILL_27_DFFSR_219 ( );
FILL FILL_28_DFFSR_219 ( );
FILL FILL_29_DFFSR_219 ( );
FILL FILL_30_DFFSR_219 ( );
FILL FILL_31_DFFSR_219 ( );
FILL FILL_32_DFFSR_219 ( );
FILL FILL_33_DFFSR_219 ( );
FILL FILL_34_DFFSR_219 ( );
FILL FILL_35_DFFSR_219 ( );
FILL FILL_36_DFFSR_219 ( );
FILL FILL_37_DFFSR_219 ( );
FILL FILL_38_DFFSR_219 ( );
FILL FILL_39_DFFSR_219 ( );
FILL FILL_40_DFFSR_219 ( );
FILL FILL_41_DFFSR_219 ( );
FILL FILL_42_DFFSR_219 ( );
FILL FILL_43_DFFSR_219 ( );
FILL FILL_44_DFFSR_219 ( );
FILL FILL_45_DFFSR_219 ( );
FILL FILL_46_DFFSR_219 ( );
FILL FILL_47_DFFSR_219 ( );
FILL FILL_48_DFFSR_219 ( );
FILL FILL_49_DFFSR_219 ( );
FILL FILL_50_DFFSR_219 ( );
FILL FILL_0_DFFSR_161 ( );
FILL FILL_1_DFFSR_161 ( );
FILL FILL_2_DFFSR_161 ( );
FILL FILL_3_DFFSR_161 ( );
FILL FILL_4_DFFSR_161 ( );
FILL FILL_5_DFFSR_161 ( );
FILL FILL_6_DFFSR_161 ( );
FILL FILL_7_DFFSR_161 ( );
FILL FILL_8_DFFSR_161 ( );
FILL FILL_9_DFFSR_161 ( );
FILL FILL_10_DFFSR_161 ( );
FILL FILL_11_DFFSR_161 ( );
FILL FILL_12_DFFSR_161 ( );
FILL FILL_13_DFFSR_161 ( );
FILL FILL_14_DFFSR_161 ( );
FILL FILL_15_DFFSR_161 ( );
FILL FILL_16_DFFSR_161 ( );
FILL FILL_17_DFFSR_161 ( );
FILL FILL_18_DFFSR_161 ( );
FILL FILL_19_DFFSR_161 ( );
FILL FILL_20_DFFSR_161 ( );
FILL FILL_21_DFFSR_161 ( );
FILL FILL_22_DFFSR_161 ( );
FILL FILL_23_DFFSR_161 ( );
FILL FILL_24_DFFSR_161 ( );
FILL FILL_25_DFFSR_161 ( );
FILL FILL_26_DFFSR_161 ( );
FILL FILL_27_DFFSR_161 ( );
FILL FILL_28_DFFSR_161 ( );
FILL FILL_29_DFFSR_161 ( );
FILL FILL_30_DFFSR_161 ( );
FILL FILL_31_DFFSR_161 ( );
FILL FILL_32_DFFSR_161 ( );
FILL FILL_33_DFFSR_161 ( );
FILL FILL_34_DFFSR_161 ( );
FILL FILL_35_DFFSR_161 ( );
FILL FILL_36_DFFSR_161 ( );
FILL FILL_37_DFFSR_161 ( );
FILL FILL_38_DFFSR_161 ( );
FILL FILL_39_DFFSR_161 ( );
FILL FILL_40_DFFSR_161 ( );
FILL FILL_41_DFFSR_161 ( );
FILL FILL_42_DFFSR_161 ( );
FILL FILL_43_DFFSR_161 ( );
FILL FILL_44_DFFSR_161 ( );
FILL FILL_45_DFFSR_161 ( );
FILL FILL_46_DFFSR_161 ( );
FILL FILL_47_DFFSR_161 ( );
FILL FILL_48_DFFSR_161 ( );
FILL FILL_49_DFFSR_161 ( );
FILL FILL_50_DFFSR_161 ( );
FILL FILL_51_DFFSR_161 ( );
FILL FILL_0_DFFSR_225 ( );
FILL FILL_1_DFFSR_225 ( );
FILL FILL_2_DFFSR_225 ( );
FILL FILL_3_DFFSR_225 ( );
FILL FILL_4_DFFSR_225 ( );
FILL FILL_5_DFFSR_225 ( );
FILL FILL_6_DFFSR_225 ( );
FILL FILL_7_DFFSR_225 ( );
FILL FILL_8_DFFSR_225 ( );
FILL FILL_9_DFFSR_225 ( );
FILL FILL_10_DFFSR_225 ( );
FILL FILL_11_DFFSR_225 ( );
FILL FILL_12_DFFSR_225 ( );
FILL FILL_13_DFFSR_225 ( );
FILL FILL_14_DFFSR_225 ( );
FILL FILL_15_DFFSR_225 ( );
FILL FILL_16_DFFSR_225 ( );
FILL FILL_17_DFFSR_225 ( );
FILL FILL_18_DFFSR_225 ( );
FILL FILL_19_DFFSR_225 ( );
FILL FILL_20_DFFSR_225 ( );
FILL FILL_21_DFFSR_225 ( );
FILL FILL_22_DFFSR_225 ( );
FILL FILL_23_DFFSR_225 ( );
FILL FILL_24_DFFSR_225 ( );
FILL FILL_25_DFFSR_225 ( );
FILL FILL_26_DFFSR_225 ( );
FILL FILL_27_DFFSR_225 ( );
FILL FILL_28_DFFSR_225 ( );
FILL FILL_29_DFFSR_225 ( );
FILL FILL_30_DFFSR_225 ( );
FILL FILL_31_DFFSR_225 ( );
FILL FILL_32_DFFSR_225 ( );
FILL FILL_33_DFFSR_225 ( );
FILL FILL_34_DFFSR_225 ( );
FILL FILL_35_DFFSR_225 ( );
FILL FILL_36_DFFSR_225 ( );
FILL FILL_37_DFFSR_225 ( );
FILL FILL_38_DFFSR_225 ( );
FILL FILL_39_DFFSR_225 ( );
FILL FILL_40_DFFSR_225 ( );
FILL FILL_41_DFFSR_225 ( );
FILL FILL_42_DFFSR_225 ( );
FILL FILL_43_DFFSR_225 ( );
FILL FILL_44_DFFSR_225 ( );
FILL FILL_45_DFFSR_225 ( );
FILL FILL_46_DFFSR_225 ( );
FILL FILL_47_DFFSR_225 ( );
FILL FILL_48_DFFSR_225 ( );
FILL FILL_49_DFFSR_225 ( );
FILL FILL_50_DFFSR_225 ( );
FILL FILL_0_DFFSR_183 ( );
FILL FILL_1_DFFSR_183 ( );
FILL FILL_2_DFFSR_183 ( );
FILL FILL_3_DFFSR_183 ( );
FILL FILL_4_DFFSR_183 ( );
FILL FILL_5_DFFSR_183 ( );
FILL FILL_6_DFFSR_183 ( );
FILL FILL_7_DFFSR_183 ( );
FILL FILL_8_DFFSR_183 ( );
FILL FILL_9_DFFSR_183 ( );
FILL FILL_10_DFFSR_183 ( );
FILL FILL_11_DFFSR_183 ( );
FILL FILL_12_DFFSR_183 ( );
FILL FILL_13_DFFSR_183 ( );
FILL FILL_14_DFFSR_183 ( );
FILL FILL_15_DFFSR_183 ( );
FILL FILL_16_DFFSR_183 ( );
FILL FILL_17_DFFSR_183 ( );
FILL FILL_18_DFFSR_183 ( );
FILL FILL_19_DFFSR_183 ( );
FILL FILL_20_DFFSR_183 ( );
FILL FILL_21_DFFSR_183 ( );
FILL FILL_22_DFFSR_183 ( );
FILL FILL_23_DFFSR_183 ( );
FILL FILL_24_DFFSR_183 ( );
FILL FILL_25_DFFSR_183 ( );
FILL FILL_26_DFFSR_183 ( );
FILL FILL_27_DFFSR_183 ( );
FILL FILL_28_DFFSR_183 ( );
FILL FILL_29_DFFSR_183 ( );
FILL FILL_30_DFFSR_183 ( );
FILL FILL_31_DFFSR_183 ( );
FILL FILL_32_DFFSR_183 ( );
FILL FILL_33_DFFSR_183 ( );
FILL FILL_34_DFFSR_183 ( );
FILL FILL_35_DFFSR_183 ( );
FILL FILL_36_DFFSR_183 ( );
FILL FILL_37_DFFSR_183 ( );
FILL FILL_38_DFFSR_183 ( );
FILL FILL_39_DFFSR_183 ( );
FILL FILL_40_DFFSR_183 ( );
FILL FILL_41_DFFSR_183 ( );
FILL FILL_42_DFFSR_183 ( );
FILL FILL_43_DFFSR_183 ( );
FILL FILL_44_DFFSR_183 ( );
FILL FILL_45_DFFSR_183 ( );
FILL FILL_46_DFFSR_183 ( );
FILL FILL_47_DFFSR_183 ( );
FILL FILL_48_DFFSR_183 ( );
FILL FILL_49_DFFSR_183 ( );
FILL FILL_50_DFFSR_183 ( );
FILL FILL_0_DFFSR_191 ( );
FILL FILL_1_DFFSR_191 ( );
FILL FILL_2_DFFSR_191 ( );
FILL FILL_3_DFFSR_191 ( );
FILL FILL_4_DFFSR_191 ( );
FILL FILL_5_DFFSR_191 ( );
FILL FILL_6_DFFSR_191 ( );
FILL FILL_7_DFFSR_191 ( );
FILL FILL_8_DFFSR_191 ( );
FILL FILL_9_DFFSR_191 ( );
FILL FILL_10_DFFSR_191 ( );
FILL FILL_11_DFFSR_191 ( );
FILL FILL_12_DFFSR_191 ( );
FILL FILL_13_DFFSR_191 ( );
FILL FILL_14_DFFSR_191 ( );
FILL FILL_15_DFFSR_191 ( );
FILL FILL_16_DFFSR_191 ( );
FILL FILL_17_DFFSR_191 ( );
FILL FILL_18_DFFSR_191 ( );
FILL FILL_19_DFFSR_191 ( );
FILL FILL_20_DFFSR_191 ( );
FILL FILL_21_DFFSR_191 ( );
FILL FILL_22_DFFSR_191 ( );
FILL FILL_23_DFFSR_191 ( );
FILL FILL_24_DFFSR_191 ( );
FILL FILL_25_DFFSR_191 ( );
FILL FILL_26_DFFSR_191 ( );
FILL FILL_27_DFFSR_191 ( );
FILL FILL_28_DFFSR_191 ( );
FILL FILL_29_DFFSR_191 ( );
FILL FILL_30_DFFSR_191 ( );
FILL FILL_31_DFFSR_191 ( );
FILL FILL_32_DFFSR_191 ( );
FILL FILL_33_DFFSR_191 ( );
FILL FILL_34_DFFSR_191 ( );
FILL FILL_35_DFFSR_191 ( );
FILL FILL_36_DFFSR_191 ( );
FILL FILL_37_DFFSR_191 ( );
FILL FILL_38_DFFSR_191 ( );
FILL FILL_39_DFFSR_191 ( );
FILL FILL_40_DFFSR_191 ( );
FILL FILL_41_DFFSR_191 ( );
FILL FILL_42_DFFSR_191 ( );
FILL FILL_43_DFFSR_191 ( );
FILL FILL_44_DFFSR_191 ( );
FILL FILL_45_DFFSR_191 ( );
FILL FILL_46_DFFSR_191 ( );
FILL FILL_47_DFFSR_191 ( );
FILL FILL_48_DFFSR_191 ( );
FILL FILL_49_DFFSR_191 ( );
FILL FILL_50_DFFSR_191 ( );
FILL FILL_51_DFFSR_191 ( );
FILL FILL_0_INVX1_137 ( );
FILL FILL_1_INVX1_137 ( );
FILL FILL_2_INVX1_137 ( );
FILL FILL_3_INVX1_137 ( );
FILL FILL_4_INVX1_137 ( );
FILL FILL_0_NAND2X1_125 ( );
FILL FILL_1_NAND2X1_125 ( );
FILL FILL_2_NAND2X1_125 ( );
FILL FILL_3_NAND2X1_125 ( );
FILL FILL_4_NAND2X1_125 ( );
FILL FILL_5_NAND2X1_125 ( );
FILL FILL_6_NAND2X1_125 ( );
FILL FILL_0_XOR2X1_2 ( );
FILL FILL_1_XOR2X1_2 ( );
FILL FILL_2_XOR2X1_2 ( );
FILL FILL_3_XOR2X1_2 ( );
FILL FILL_4_XOR2X1_2 ( );
FILL FILL_5_XOR2X1_2 ( );
FILL FILL_6_XOR2X1_2 ( );
FILL FILL_7_XOR2X1_2 ( );
FILL FILL_8_XOR2X1_2 ( );
FILL FILL_9_XOR2X1_2 ( );
FILL FILL_10_XOR2X1_2 ( );
FILL FILL_11_XOR2X1_2 ( );
FILL FILL_12_XOR2X1_2 ( );
FILL FILL_13_XOR2X1_2 ( );
FILL FILL_14_XOR2X1_2 ( );
FILL FILL_15_XOR2X1_2 ( );
FILL FILL_0_OAI21X1_26 ( );
FILL FILL_1_OAI21X1_26 ( );
FILL FILL_2_OAI21X1_26 ( );
FILL FILL_3_OAI21X1_26 ( );
FILL FILL_4_OAI21X1_26 ( );
FILL FILL_5_OAI21X1_26 ( );
FILL FILL_6_OAI21X1_26 ( );
FILL FILL_7_OAI21X1_26 ( );
FILL FILL_8_OAI21X1_26 ( );
FILL FILL_9_OAI21X1_26 ( );
FILL FILL_0_OAI21X1_93 ( );
FILL FILL_1_OAI21X1_93 ( );
FILL FILL_2_OAI21X1_93 ( );
FILL FILL_3_OAI21X1_93 ( );
FILL FILL_4_OAI21X1_93 ( );
FILL FILL_5_OAI21X1_93 ( );
FILL FILL_6_OAI21X1_93 ( );
FILL FILL_7_OAI21X1_93 ( );
FILL FILL_8_OAI21X1_93 ( );
FILL FILL_9_OAI21X1_93 ( );
FILL FILL_0_INVX1_155 ( );
FILL FILL_1_INVX1_155 ( );
FILL FILL_2_INVX1_155 ( );
FILL FILL_3_INVX1_155 ( );
FILL FILL_4_INVX1_155 ( );
FILL FILL_0_AOI21X1_18 ( );
FILL FILL_1_AOI21X1_18 ( );
FILL FILL_2_AOI21X1_18 ( );
FILL FILL_3_AOI21X1_18 ( );
FILL FILL_4_AOI21X1_18 ( );
FILL FILL_5_AOI21X1_18 ( );
FILL FILL_6_AOI21X1_18 ( );
FILL FILL_7_AOI21X1_18 ( );
FILL FILL_8_AOI21X1_18 ( );
FILL FILL_0_INVX1_140 ( );
FILL FILL_1_INVX1_140 ( );
FILL FILL_2_INVX1_140 ( );
FILL FILL_3_INVX1_140 ( );
FILL FILL_0_OAI21X1_29 ( );
FILL FILL_1_OAI21X1_29 ( );
FILL FILL_2_OAI21X1_29 ( );
FILL FILL_3_OAI21X1_29 ( );
FILL FILL_4_OAI21X1_29 ( );
FILL FILL_5_OAI21X1_29 ( );
FILL FILL_6_OAI21X1_29 ( );
FILL FILL_7_OAI21X1_29 ( );
FILL FILL_8_OAI21X1_29 ( );
FILL FILL_0_AOI21X1_7 ( );
FILL FILL_1_AOI21X1_7 ( );
FILL FILL_2_AOI21X1_7 ( );
FILL FILL_3_AOI21X1_7 ( );
FILL FILL_4_AOI21X1_7 ( );
FILL FILL_5_AOI21X1_7 ( );
FILL FILL_6_AOI21X1_7 ( );
FILL FILL_7_AOI21X1_7 ( );
FILL FILL_8_AOI21X1_7 ( );
FILL FILL_9_AOI21X1_7 ( );
FILL FILL_0_NOR2X1_68 ( );
FILL FILL_1_NOR2X1_68 ( );
FILL FILL_2_NOR2X1_68 ( );
FILL FILL_3_NOR2X1_68 ( );
FILL FILL_4_NOR2X1_68 ( );
FILL FILL_5_NOR2X1_68 ( );
FILL FILL_6_NOR2X1_68 ( );
FILL FILL_0_AND2X2_30 ( );
FILL FILL_1_AND2X2_30 ( );
FILL FILL_2_AND2X2_30 ( );
FILL FILL_3_AND2X2_30 ( );
FILL FILL_4_AND2X2_30 ( );
FILL FILL_5_AND2X2_30 ( );
FILL FILL_6_AND2X2_30 ( );
FILL FILL_7_AND2X2_30 ( );
FILL FILL_8_AND2X2_30 ( );
FILL FILL_0_NAND2X1_126 ( );
FILL FILL_1_NAND2X1_126 ( );
FILL FILL_2_NAND2X1_126 ( );
FILL FILL_3_NAND2X1_126 ( );
FILL FILL_4_NAND2X1_126 ( );
FILL FILL_5_NAND2X1_126 ( );
FILL FILL_6_NAND2X1_126 ( );
FILL FILL_0_BUFX2_36 ( );
FILL FILL_1_BUFX2_36 ( );
FILL FILL_2_BUFX2_36 ( );
FILL FILL_3_BUFX2_36 ( );
FILL FILL_4_BUFX2_36 ( );
FILL FILL_5_BUFX2_36 ( );
FILL FILL_6_BUFX2_36 ( );
FILL FILL_0_AOI21X1_58 ( );
FILL FILL_1_AOI21X1_58 ( );
FILL FILL_2_AOI21X1_58 ( );
FILL FILL_3_AOI21X1_58 ( );
FILL FILL_4_AOI21X1_58 ( );
FILL FILL_5_AOI21X1_58 ( );
FILL FILL_6_AOI21X1_58 ( );
FILL FILL_7_AOI21X1_58 ( );
FILL FILL_8_AOI21X1_58 ( );
FILL FILL_0_DFFPOSX1_36 ( );
FILL FILL_1_DFFPOSX1_36 ( );
FILL FILL_2_DFFPOSX1_36 ( );
FILL FILL_3_DFFPOSX1_36 ( );
FILL FILL_4_DFFPOSX1_36 ( );
FILL FILL_5_DFFPOSX1_36 ( );
FILL FILL_6_DFFPOSX1_36 ( );
FILL FILL_7_DFFPOSX1_36 ( );
FILL FILL_8_DFFPOSX1_36 ( );
FILL FILL_9_DFFPOSX1_36 ( );
FILL FILL_10_DFFPOSX1_36 ( );
FILL FILL_11_DFFPOSX1_36 ( );
FILL FILL_12_DFFPOSX1_36 ( );
FILL FILL_13_DFFPOSX1_36 ( );
FILL FILL_14_DFFPOSX1_36 ( );
FILL FILL_15_DFFPOSX1_36 ( );
FILL FILL_16_DFFPOSX1_36 ( );
FILL FILL_17_DFFPOSX1_36 ( );
FILL FILL_18_DFFPOSX1_36 ( );
FILL FILL_19_DFFPOSX1_36 ( );
FILL FILL_20_DFFPOSX1_36 ( );
FILL FILL_21_DFFPOSX1_36 ( );
FILL FILL_22_DFFPOSX1_36 ( );
FILL FILL_23_DFFPOSX1_36 ( );
FILL FILL_24_DFFPOSX1_36 ( );
FILL FILL_25_DFFPOSX1_36 ( );
FILL FILL_26_DFFPOSX1_36 ( );
FILL FILL_27_DFFPOSX1_36 ( );
FILL FILL_0_DFFSR_212 ( );
FILL FILL_1_DFFSR_212 ( );
FILL FILL_2_DFFSR_212 ( );
FILL FILL_3_DFFSR_212 ( );
FILL FILL_4_DFFSR_212 ( );
FILL FILL_5_DFFSR_212 ( );
FILL FILL_6_DFFSR_212 ( );
FILL FILL_7_DFFSR_212 ( );
FILL FILL_8_DFFSR_212 ( );
FILL FILL_9_DFFSR_212 ( );
FILL FILL_10_DFFSR_212 ( );
FILL FILL_11_DFFSR_212 ( );
FILL FILL_12_DFFSR_212 ( );
FILL FILL_13_DFFSR_212 ( );
FILL FILL_14_DFFSR_212 ( );
FILL FILL_15_DFFSR_212 ( );
FILL FILL_16_DFFSR_212 ( );
FILL FILL_17_DFFSR_212 ( );
FILL FILL_18_DFFSR_212 ( );
FILL FILL_19_DFFSR_212 ( );
FILL FILL_20_DFFSR_212 ( );
FILL FILL_21_DFFSR_212 ( );
FILL FILL_22_DFFSR_212 ( );
FILL FILL_23_DFFSR_212 ( );
FILL FILL_24_DFFSR_212 ( );
FILL FILL_25_DFFSR_212 ( );
FILL FILL_26_DFFSR_212 ( );
FILL FILL_27_DFFSR_212 ( );
FILL FILL_28_DFFSR_212 ( );
FILL FILL_29_DFFSR_212 ( );
FILL FILL_30_DFFSR_212 ( );
FILL FILL_31_DFFSR_212 ( );
FILL FILL_32_DFFSR_212 ( );
FILL FILL_33_DFFSR_212 ( );
FILL FILL_34_DFFSR_212 ( );
FILL FILL_35_DFFSR_212 ( );
FILL FILL_36_DFFSR_212 ( );
FILL FILL_37_DFFSR_212 ( );
FILL FILL_38_DFFSR_212 ( );
FILL FILL_39_DFFSR_212 ( );
FILL FILL_40_DFFSR_212 ( );
FILL FILL_41_DFFSR_212 ( );
FILL FILL_42_DFFSR_212 ( );
FILL FILL_43_DFFSR_212 ( );
FILL FILL_44_DFFSR_212 ( );
FILL FILL_45_DFFSR_212 ( );
FILL FILL_46_DFFSR_212 ( );
FILL FILL_47_DFFSR_212 ( );
FILL FILL_48_DFFSR_212 ( );
FILL FILL_49_DFFSR_212 ( );
FILL FILL_50_DFFSR_212 ( );
FILL FILL_0_DFFSR_206 ( );
FILL FILL_1_DFFSR_206 ( );
FILL FILL_2_DFFSR_206 ( );
FILL FILL_3_DFFSR_206 ( );
FILL FILL_4_DFFSR_206 ( );
FILL FILL_5_DFFSR_206 ( );
FILL FILL_6_DFFSR_206 ( );
FILL FILL_7_DFFSR_206 ( );
FILL FILL_8_DFFSR_206 ( );
FILL FILL_9_DFFSR_206 ( );
FILL FILL_10_DFFSR_206 ( );
FILL FILL_11_DFFSR_206 ( );
FILL FILL_12_DFFSR_206 ( );
FILL FILL_13_DFFSR_206 ( );
FILL FILL_14_DFFSR_206 ( );
FILL FILL_15_DFFSR_206 ( );
FILL FILL_16_DFFSR_206 ( );
FILL FILL_17_DFFSR_206 ( );
FILL FILL_18_DFFSR_206 ( );
FILL FILL_19_DFFSR_206 ( );
FILL FILL_20_DFFSR_206 ( );
FILL FILL_21_DFFSR_206 ( );
FILL FILL_22_DFFSR_206 ( );
FILL FILL_23_DFFSR_206 ( );
FILL FILL_24_DFFSR_206 ( );
FILL FILL_25_DFFSR_206 ( );
FILL FILL_26_DFFSR_206 ( );
FILL FILL_27_DFFSR_206 ( );
FILL FILL_28_DFFSR_206 ( );
FILL FILL_29_DFFSR_206 ( );
FILL FILL_30_DFFSR_206 ( );
FILL FILL_31_DFFSR_206 ( );
FILL FILL_32_DFFSR_206 ( );
FILL FILL_33_DFFSR_206 ( );
FILL FILL_34_DFFSR_206 ( );
FILL FILL_35_DFFSR_206 ( );
FILL FILL_36_DFFSR_206 ( );
FILL FILL_37_DFFSR_206 ( );
FILL FILL_38_DFFSR_206 ( );
FILL FILL_39_DFFSR_206 ( );
FILL FILL_40_DFFSR_206 ( );
FILL FILL_41_DFFSR_206 ( );
FILL FILL_42_DFFSR_206 ( );
FILL FILL_43_DFFSR_206 ( );
FILL FILL_44_DFFSR_206 ( );
FILL FILL_45_DFFSR_206 ( );
FILL FILL_46_DFFSR_206 ( );
FILL FILL_47_DFFSR_206 ( );
FILL FILL_48_DFFSR_206 ( );
FILL FILL_49_DFFSR_206 ( );
FILL FILL_50_DFFSR_206 ( );
FILL FILL_0_INVX1_100 ( );
FILL FILL_1_INVX1_100 ( );
FILL FILL_2_INVX1_100 ( );
FILL FILL_3_INVX1_100 ( );
FILL FILL_0_INVX1_87 ( );
FILL FILL_1_INVX1_87 ( );
FILL FILL_2_INVX1_87 ( );
FILL FILL_3_INVX1_87 ( );
FILL FILL_0_DFFSR_156 ( );
FILL FILL_1_DFFSR_156 ( );
FILL FILL_2_DFFSR_156 ( );
FILL FILL_3_DFFSR_156 ( );
FILL FILL_4_DFFSR_156 ( );
FILL FILL_5_DFFSR_156 ( );
FILL FILL_6_DFFSR_156 ( );
FILL FILL_7_DFFSR_156 ( );
FILL FILL_8_DFFSR_156 ( );
FILL FILL_9_DFFSR_156 ( );
FILL FILL_10_DFFSR_156 ( );
FILL FILL_11_DFFSR_156 ( );
FILL FILL_12_DFFSR_156 ( );
FILL FILL_13_DFFSR_156 ( );
FILL FILL_14_DFFSR_156 ( );
FILL FILL_15_DFFSR_156 ( );
FILL FILL_16_DFFSR_156 ( );
FILL FILL_17_DFFSR_156 ( );
FILL FILL_18_DFFSR_156 ( );
FILL FILL_19_DFFSR_156 ( );
FILL FILL_20_DFFSR_156 ( );
FILL FILL_21_DFFSR_156 ( );
FILL FILL_22_DFFSR_156 ( );
FILL FILL_23_DFFSR_156 ( );
FILL FILL_24_DFFSR_156 ( );
FILL FILL_25_DFFSR_156 ( );
FILL FILL_26_DFFSR_156 ( );
FILL FILL_27_DFFSR_156 ( );
FILL FILL_28_DFFSR_156 ( );
FILL FILL_29_DFFSR_156 ( );
FILL FILL_30_DFFSR_156 ( );
FILL FILL_31_DFFSR_156 ( );
FILL FILL_32_DFFSR_156 ( );
FILL FILL_33_DFFSR_156 ( );
FILL FILL_34_DFFSR_156 ( );
FILL FILL_35_DFFSR_156 ( );
FILL FILL_36_DFFSR_156 ( );
FILL FILL_37_DFFSR_156 ( );
FILL FILL_38_DFFSR_156 ( );
FILL FILL_39_DFFSR_156 ( );
FILL FILL_40_DFFSR_156 ( );
FILL FILL_41_DFFSR_156 ( );
FILL FILL_42_DFFSR_156 ( );
FILL FILL_43_DFFSR_156 ( );
FILL FILL_44_DFFSR_156 ( );
FILL FILL_45_DFFSR_156 ( );
FILL FILL_46_DFFSR_156 ( );
FILL FILL_47_DFFSR_156 ( );
FILL FILL_48_DFFSR_156 ( );
FILL FILL_49_DFFSR_156 ( );
FILL FILL_50_DFFSR_156 ( );
FILL FILL_0_BUFX2_90 ( );
FILL FILL_1_BUFX2_90 ( );
FILL FILL_2_BUFX2_90 ( );
FILL FILL_3_BUFX2_90 ( );
FILL FILL_4_BUFX2_90 ( );
FILL FILL_5_BUFX2_90 ( );
FILL FILL_6_BUFX2_90 ( );
FILL FILL_0_DFFSR_233 ( );
FILL FILL_1_DFFSR_233 ( );
FILL FILL_2_DFFSR_233 ( );
FILL FILL_3_DFFSR_233 ( );
FILL FILL_4_DFFSR_233 ( );
FILL FILL_5_DFFSR_233 ( );
FILL FILL_6_DFFSR_233 ( );
FILL FILL_7_DFFSR_233 ( );
FILL FILL_8_DFFSR_233 ( );
FILL FILL_9_DFFSR_233 ( );
FILL FILL_10_DFFSR_233 ( );
FILL FILL_11_DFFSR_233 ( );
FILL FILL_12_DFFSR_233 ( );
FILL FILL_13_DFFSR_233 ( );
FILL FILL_14_DFFSR_233 ( );
FILL FILL_15_DFFSR_233 ( );
FILL FILL_16_DFFSR_233 ( );
FILL FILL_17_DFFSR_233 ( );
FILL FILL_18_DFFSR_233 ( );
FILL FILL_19_DFFSR_233 ( );
FILL FILL_20_DFFSR_233 ( );
FILL FILL_21_DFFSR_233 ( );
FILL FILL_22_DFFSR_233 ( );
FILL FILL_23_DFFSR_233 ( );
FILL FILL_24_DFFSR_233 ( );
FILL FILL_25_DFFSR_233 ( );
FILL FILL_26_DFFSR_233 ( );
FILL FILL_27_DFFSR_233 ( );
FILL FILL_28_DFFSR_233 ( );
FILL FILL_29_DFFSR_233 ( );
FILL FILL_30_DFFSR_233 ( );
FILL FILL_31_DFFSR_233 ( );
FILL FILL_32_DFFSR_233 ( );
FILL FILL_33_DFFSR_233 ( );
FILL FILL_34_DFFSR_233 ( );
FILL FILL_35_DFFSR_233 ( );
FILL FILL_36_DFFSR_233 ( );
FILL FILL_37_DFFSR_233 ( );
FILL FILL_38_DFFSR_233 ( );
FILL FILL_39_DFFSR_233 ( );
FILL FILL_40_DFFSR_233 ( );
FILL FILL_41_DFFSR_233 ( );
FILL FILL_42_DFFSR_233 ( );
FILL FILL_43_DFFSR_233 ( );
FILL FILL_44_DFFSR_233 ( );
FILL FILL_45_DFFSR_233 ( );
FILL FILL_46_DFFSR_233 ( );
FILL FILL_47_DFFSR_233 ( );
FILL FILL_48_DFFSR_233 ( );
FILL FILL_49_DFFSR_233 ( );
FILL FILL_50_DFFSR_233 ( );
FILL FILL_0_DFFSR_193 ( );
FILL FILL_1_DFFSR_193 ( );
FILL FILL_2_DFFSR_193 ( );
FILL FILL_3_DFFSR_193 ( );
FILL FILL_4_DFFSR_193 ( );
FILL FILL_5_DFFSR_193 ( );
FILL FILL_6_DFFSR_193 ( );
FILL FILL_7_DFFSR_193 ( );
FILL FILL_8_DFFSR_193 ( );
FILL FILL_9_DFFSR_193 ( );
FILL FILL_10_DFFSR_193 ( );
FILL FILL_11_DFFSR_193 ( );
FILL FILL_12_DFFSR_193 ( );
FILL FILL_13_DFFSR_193 ( );
FILL FILL_14_DFFSR_193 ( );
FILL FILL_15_DFFSR_193 ( );
FILL FILL_16_DFFSR_193 ( );
FILL FILL_17_DFFSR_193 ( );
FILL FILL_18_DFFSR_193 ( );
FILL FILL_19_DFFSR_193 ( );
FILL FILL_20_DFFSR_193 ( );
FILL FILL_21_DFFSR_193 ( );
FILL FILL_22_DFFSR_193 ( );
FILL FILL_23_DFFSR_193 ( );
FILL FILL_24_DFFSR_193 ( );
FILL FILL_25_DFFSR_193 ( );
FILL FILL_26_DFFSR_193 ( );
FILL FILL_27_DFFSR_193 ( );
FILL FILL_28_DFFSR_193 ( );
FILL FILL_29_DFFSR_193 ( );
FILL FILL_30_DFFSR_193 ( );
FILL FILL_31_DFFSR_193 ( );
FILL FILL_32_DFFSR_193 ( );
FILL FILL_33_DFFSR_193 ( );
FILL FILL_34_DFFSR_193 ( );
FILL FILL_35_DFFSR_193 ( );
FILL FILL_36_DFFSR_193 ( );
FILL FILL_37_DFFSR_193 ( );
FILL FILL_38_DFFSR_193 ( );
FILL FILL_39_DFFSR_193 ( );
FILL FILL_40_DFFSR_193 ( );
FILL FILL_41_DFFSR_193 ( );
FILL FILL_42_DFFSR_193 ( );
FILL FILL_43_DFFSR_193 ( );
FILL FILL_44_DFFSR_193 ( );
FILL FILL_45_DFFSR_193 ( );
FILL FILL_46_DFFSR_193 ( );
FILL FILL_47_DFFSR_193 ( );
FILL FILL_48_DFFSR_193 ( );
FILL FILL_49_DFFSR_193 ( );
FILL FILL_50_DFFSR_193 ( );
FILL FILL_0_DFFSR_175 ( );
FILL FILL_1_DFFSR_175 ( );
FILL FILL_2_DFFSR_175 ( );
FILL FILL_3_DFFSR_175 ( );
FILL FILL_4_DFFSR_175 ( );
FILL FILL_5_DFFSR_175 ( );
FILL FILL_6_DFFSR_175 ( );
FILL FILL_7_DFFSR_175 ( );
FILL FILL_8_DFFSR_175 ( );
FILL FILL_9_DFFSR_175 ( );
FILL FILL_10_DFFSR_175 ( );
FILL FILL_11_DFFSR_175 ( );
FILL FILL_12_DFFSR_175 ( );
FILL FILL_13_DFFSR_175 ( );
FILL FILL_14_DFFSR_175 ( );
FILL FILL_15_DFFSR_175 ( );
FILL FILL_16_DFFSR_175 ( );
FILL FILL_17_DFFSR_175 ( );
FILL FILL_18_DFFSR_175 ( );
FILL FILL_19_DFFSR_175 ( );
FILL FILL_20_DFFSR_175 ( );
FILL FILL_21_DFFSR_175 ( );
FILL FILL_22_DFFSR_175 ( );
FILL FILL_23_DFFSR_175 ( );
FILL FILL_24_DFFSR_175 ( );
FILL FILL_25_DFFSR_175 ( );
FILL FILL_26_DFFSR_175 ( );
FILL FILL_27_DFFSR_175 ( );
FILL FILL_28_DFFSR_175 ( );
FILL FILL_29_DFFSR_175 ( );
FILL FILL_30_DFFSR_175 ( );
FILL FILL_31_DFFSR_175 ( );
FILL FILL_32_DFFSR_175 ( );
FILL FILL_33_DFFSR_175 ( );
FILL FILL_34_DFFSR_175 ( );
FILL FILL_35_DFFSR_175 ( );
FILL FILL_36_DFFSR_175 ( );
FILL FILL_37_DFFSR_175 ( );
FILL FILL_38_DFFSR_175 ( );
FILL FILL_39_DFFSR_175 ( );
FILL FILL_40_DFFSR_175 ( );
FILL FILL_41_DFFSR_175 ( );
FILL FILL_42_DFFSR_175 ( );
FILL FILL_43_DFFSR_175 ( );
FILL FILL_44_DFFSR_175 ( );
FILL FILL_45_DFFSR_175 ( );
FILL FILL_46_DFFSR_175 ( );
FILL FILL_47_DFFSR_175 ( );
FILL FILL_48_DFFSR_175 ( );
FILL FILL_49_DFFSR_175 ( );
FILL FILL_50_DFFSR_175 ( );
FILL FILL_0_BUFX2_76 ( );
FILL FILL_1_BUFX2_76 ( );
FILL FILL_2_BUFX2_76 ( );
FILL FILL_3_BUFX2_76 ( );
FILL FILL_4_BUFX2_76 ( );
FILL FILL_5_BUFX2_76 ( );
FILL FILL_6_BUFX2_76 ( );
FILL FILL_0_NAND3X1_192 ( );
FILL FILL_1_NAND3X1_192 ( );
FILL FILL_2_NAND3X1_192 ( );
FILL FILL_3_NAND3X1_192 ( );
FILL FILL_4_NAND3X1_192 ( );
FILL FILL_5_NAND3X1_192 ( );
FILL FILL_6_NAND3X1_192 ( );
FILL FILL_7_NAND3X1_192 ( );
FILL FILL_8_NAND3X1_192 ( );
FILL FILL_0_OR2X2_2 ( );
FILL FILL_1_OR2X2_2 ( );
FILL FILL_2_OR2X2_2 ( );
FILL FILL_3_OR2X2_2 ( );
FILL FILL_4_OR2X2_2 ( );
FILL FILL_5_OR2X2_2 ( );
FILL FILL_6_OR2X2_2 ( );
FILL FILL_7_OR2X2_2 ( );
FILL FILL_8_OR2X2_2 ( );
FILL FILL_9_OR2X2_2 ( );
FILL FILL_0_NAND2X1_61 ( );
FILL FILL_1_NAND2X1_61 ( );
FILL FILL_2_NAND2X1_61 ( );
FILL FILL_3_NAND2X1_61 ( );
FILL FILL_4_NAND2X1_61 ( );
FILL FILL_5_NAND2X1_61 ( );
FILL FILL_6_NAND2X1_61 ( );
FILL FILL_0_INVX1_136 ( );
FILL FILL_1_INVX1_136 ( );
FILL FILL_2_INVX1_136 ( );
FILL FILL_3_INVX1_136 ( );
FILL FILL_0_NAND2X1_124 ( );
FILL FILL_1_NAND2X1_124 ( );
FILL FILL_2_NAND2X1_124 ( );
FILL FILL_3_NAND2X1_124 ( );
FILL FILL_4_NAND2X1_124 ( );
FILL FILL_5_NAND2X1_124 ( );
FILL FILL_6_NAND2X1_124 ( );
FILL FILL_0_INVX1_190 ( );
FILL FILL_1_INVX1_190 ( );
FILL FILL_2_INVX1_190 ( );
FILL FILL_3_INVX1_190 ( );
FILL FILL_0_NAND2X1_70 ( );
FILL FILL_1_NAND2X1_70 ( );
FILL FILL_2_NAND2X1_70 ( );
FILL FILL_3_NAND2X1_70 ( );
FILL FILL_4_NAND2X1_70 ( );
FILL FILL_5_NAND2X1_70 ( );
FILL FILL_6_NAND2X1_70 ( );
FILL FILL_0_XOR2X1_3 ( );
FILL FILL_1_XOR2X1_3 ( );
FILL FILL_2_XOR2X1_3 ( );
FILL FILL_3_XOR2X1_3 ( );
FILL FILL_4_XOR2X1_3 ( );
FILL FILL_5_XOR2X1_3 ( );
FILL FILL_6_XOR2X1_3 ( );
FILL FILL_7_XOR2X1_3 ( );
FILL FILL_8_XOR2X1_3 ( );
FILL FILL_9_XOR2X1_3 ( );
FILL FILL_10_XOR2X1_3 ( );
FILL FILL_11_XOR2X1_3 ( );
FILL FILL_12_XOR2X1_3 ( );
FILL FILL_13_XOR2X1_3 ( );
FILL FILL_14_XOR2X1_3 ( );
FILL FILL_15_XOR2X1_3 ( );
FILL FILL_16_XOR2X1_3 ( );
FILL FILL_0_DFFPOSX1_44 ( );
FILL FILL_1_DFFPOSX1_44 ( );
FILL FILL_2_DFFPOSX1_44 ( );
FILL FILL_3_DFFPOSX1_44 ( );
FILL FILL_4_DFFPOSX1_44 ( );
FILL FILL_5_DFFPOSX1_44 ( );
FILL FILL_6_DFFPOSX1_44 ( );
FILL FILL_7_DFFPOSX1_44 ( );
FILL FILL_8_DFFPOSX1_44 ( );
FILL FILL_9_DFFPOSX1_44 ( );
FILL FILL_10_DFFPOSX1_44 ( );
FILL FILL_11_DFFPOSX1_44 ( );
FILL FILL_12_DFFPOSX1_44 ( );
FILL FILL_13_DFFPOSX1_44 ( );
FILL FILL_14_DFFPOSX1_44 ( );
FILL FILL_15_DFFPOSX1_44 ( );
FILL FILL_16_DFFPOSX1_44 ( );
FILL FILL_17_DFFPOSX1_44 ( );
FILL FILL_18_DFFPOSX1_44 ( );
FILL FILL_19_DFFPOSX1_44 ( );
FILL FILL_20_DFFPOSX1_44 ( );
FILL FILL_21_DFFPOSX1_44 ( );
FILL FILL_22_DFFPOSX1_44 ( );
FILL FILL_23_DFFPOSX1_44 ( );
FILL FILL_24_DFFPOSX1_44 ( );
FILL FILL_25_DFFPOSX1_44 ( );
FILL FILL_26_DFFPOSX1_44 ( );
FILL FILL_27_DFFPOSX1_44 ( );
FILL FILL_0_OAI21X1_27 ( );
FILL FILL_1_OAI21X1_27 ( );
FILL FILL_2_OAI21X1_27 ( );
FILL FILL_3_OAI21X1_27 ( );
FILL FILL_4_OAI21X1_27 ( );
FILL FILL_5_OAI21X1_27 ( );
FILL FILL_6_OAI21X1_27 ( );
FILL FILL_7_OAI21X1_27 ( );
FILL FILL_8_OAI21X1_27 ( );
FILL FILL_0_DFFPOSX1_5 ( );
FILL FILL_1_DFFPOSX1_5 ( );
FILL FILL_2_DFFPOSX1_5 ( );
FILL FILL_3_DFFPOSX1_5 ( );
FILL FILL_4_DFFPOSX1_5 ( );
FILL FILL_5_DFFPOSX1_5 ( );
FILL FILL_6_DFFPOSX1_5 ( );
FILL FILL_7_DFFPOSX1_5 ( );
FILL FILL_8_DFFPOSX1_5 ( );
FILL FILL_9_DFFPOSX1_5 ( );
FILL FILL_10_DFFPOSX1_5 ( );
FILL FILL_11_DFFPOSX1_5 ( );
FILL FILL_12_DFFPOSX1_5 ( );
FILL FILL_13_DFFPOSX1_5 ( );
FILL FILL_14_DFFPOSX1_5 ( );
FILL FILL_15_DFFPOSX1_5 ( );
FILL FILL_16_DFFPOSX1_5 ( );
FILL FILL_17_DFFPOSX1_5 ( );
FILL FILL_18_DFFPOSX1_5 ( );
FILL FILL_19_DFFPOSX1_5 ( );
FILL FILL_20_DFFPOSX1_5 ( );
FILL FILL_21_DFFPOSX1_5 ( );
FILL FILL_22_DFFPOSX1_5 ( );
FILL FILL_23_DFFPOSX1_5 ( );
FILL FILL_24_DFFPOSX1_5 ( );
FILL FILL_25_DFFPOSX1_5 ( );
FILL FILL_26_DFFPOSX1_5 ( );
FILL FILL_27_DFFPOSX1_5 ( );
FILL FILL_0_NAND2X1_147 ( );
FILL FILL_1_NAND2X1_147 ( );
FILL FILL_2_NAND2X1_147 ( );
FILL FILL_3_NAND2X1_147 ( );
FILL FILL_4_NAND2X1_147 ( );
FILL FILL_5_NAND2X1_147 ( );
FILL FILL_6_NAND2X1_147 ( );
FILL FILL_0_DFFPOSX1_34 ( );
FILL FILL_1_DFFPOSX1_34 ( );
FILL FILL_2_DFFPOSX1_34 ( );
FILL FILL_3_DFFPOSX1_34 ( );
FILL FILL_4_DFFPOSX1_34 ( );
FILL FILL_5_DFFPOSX1_34 ( );
FILL FILL_6_DFFPOSX1_34 ( );
FILL FILL_7_DFFPOSX1_34 ( );
FILL FILL_8_DFFPOSX1_34 ( );
FILL FILL_9_DFFPOSX1_34 ( );
FILL FILL_10_DFFPOSX1_34 ( );
FILL FILL_11_DFFPOSX1_34 ( );
FILL FILL_12_DFFPOSX1_34 ( );
FILL FILL_13_DFFPOSX1_34 ( );
FILL FILL_14_DFFPOSX1_34 ( );
FILL FILL_15_DFFPOSX1_34 ( );
FILL FILL_16_DFFPOSX1_34 ( );
FILL FILL_17_DFFPOSX1_34 ( );
FILL FILL_18_DFFPOSX1_34 ( );
FILL FILL_19_DFFPOSX1_34 ( );
FILL FILL_20_DFFPOSX1_34 ( );
FILL FILL_21_DFFPOSX1_34 ( );
FILL FILL_22_DFFPOSX1_34 ( );
FILL FILL_23_DFFPOSX1_34 ( );
FILL FILL_24_DFFPOSX1_34 ( );
FILL FILL_25_DFFPOSX1_34 ( );
FILL FILL_26_DFFPOSX1_34 ( );
FILL FILL_27_DFFPOSX1_34 ( );
FILL FILL_0_NAND2X1_149 ( );
FILL FILL_1_NAND2X1_149 ( );
FILL FILL_2_NAND2X1_149 ( );
FILL FILL_3_NAND2X1_149 ( );
FILL FILL_4_NAND2X1_149 ( );
FILL FILL_5_NAND2X1_149 ( );
FILL FILL_6_NAND2X1_149 ( );
FILL FILL_0_DFFPOSX1_43 ( );
FILL FILL_1_DFFPOSX1_43 ( );
FILL FILL_2_DFFPOSX1_43 ( );
FILL FILL_3_DFFPOSX1_43 ( );
FILL FILL_4_DFFPOSX1_43 ( );
FILL FILL_5_DFFPOSX1_43 ( );
FILL FILL_6_DFFPOSX1_43 ( );
FILL FILL_7_DFFPOSX1_43 ( );
FILL FILL_8_DFFPOSX1_43 ( );
FILL FILL_9_DFFPOSX1_43 ( );
FILL FILL_10_DFFPOSX1_43 ( );
FILL FILL_11_DFFPOSX1_43 ( );
FILL FILL_12_DFFPOSX1_43 ( );
FILL FILL_13_DFFPOSX1_43 ( );
FILL FILL_14_DFFPOSX1_43 ( );
FILL FILL_15_DFFPOSX1_43 ( );
FILL FILL_16_DFFPOSX1_43 ( );
FILL FILL_17_DFFPOSX1_43 ( );
FILL FILL_18_DFFPOSX1_43 ( );
FILL FILL_19_DFFPOSX1_43 ( );
FILL FILL_20_DFFPOSX1_43 ( );
FILL FILL_21_DFFPOSX1_43 ( );
FILL FILL_22_DFFPOSX1_43 ( );
FILL FILL_23_DFFPOSX1_43 ( );
FILL FILL_24_DFFPOSX1_43 ( );
FILL FILL_25_DFFPOSX1_43 ( );
FILL FILL_26_DFFPOSX1_43 ( );
FILL FILL_27_DFFPOSX1_43 ( );
FILL FILL_0_DFFSR_164 ( );
FILL FILL_1_DFFSR_164 ( );
FILL FILL_2_DFFSR_164 ( );
FILL FILL_3_DFFSR_164 ( );
FILL FILL_4_DFFSR_164 ( );
FILL FILL_5_DFFSR_164 ( );
FILL FILL_6_DFFSR_164 ( );
FILL FILL_7_DFFSR_164 ( );
FILL FILL_8_DFFSR_164 ( );
FILL FILL_9_DFFSR_164 ( );
FILL FILL_10_DFFSR_164 ( );
FILL FILL_11_DFFSR_164 ( );
FILL FILL_12_DFFSR_164 ( );
FILL FILL_13_DFFSR_164 ( );
FILL FILL_14_DFFSR_164 ( );
FILL FILL_15_DFFSR_164 ( );
FILL FILL_16_DFFSR_164 ( );
FILL FILL_17_DFFSR_164 ( );
FILL FILL_18_DFFSR_164 ( );
FILL FILL_19_DFFSR_164 ( );
FILL FILL_20_DFFSR_164 ( );
FILL FILL_21_DFFSR_164 ( );
FILL FILL_22_DFFSR_164 ( );
FILL FILL_23_DFFSR_164 ( );
FILL FILL_24_DFFSR_164 ( );
FILL FILL_25_DFFSR_164 ( );
FILL FILL_26_DFFSR_164 ( );
FILL FILL_27_DFFSR_164 ( );
FILL FILL_28_DFFSR_164 ( );
FILL FILL_29_DFFSR_164 ( );
FILL FILL_30_DFFSR_164 ( );
FILL FILL_31_DFFSR_164 ( );
FILL FILL_32_DFFSR_164 ( );
FILL FILL_33_DFFSR_164 ( );
FILL FILL_34_DFFSR_164 ( );
FILL FILL_35_DFFSR_164 ( );
FILL FILL_36_DFFSR_164 ( );
FILL FILL_37_DFFSR_164 ( );
FILL FILL_38_DFFSR_164 ( );
FILL FILL_39_DFFSR_164 ( );
FILL FILL_40_DFFSR_164 ( );
FILL FILL_41_DFFSR_164 ( );
FILL FILL_42_DFFSR_164 ( );
FILL FILL_43_DFFSR_164 ( );
FILL FILL_44_DFFSR_164 ( );
FILL FILL_45_DFFSR_164 ( );
FILL FILL_46_DFFSR_164 ( );
FILL FILL_47_DFFSR_164 ( );
FILL FILL_48_DFFSR_164 ( );
FILL FILL_49_DFFSR_164 ( );
FILL FILL_50_DFFSR_164 ( );
FILL FILL_51_DFFSR_164 ( );
FILL FILL_0_BUFX2_60 ( );
FILL FILL_1_BUFX2_60 ( );
FILL FILL_2_BUFX2_60 ( );
FILL FILL_3_BUFX2_60 ( );
FILL FILL_4_BUFX2_60 ( );
FILL FILL_5_BUFX2_60 ( );
FILL FILL_6_BUFX2_60 ( );
FILL FILL_0_AOI22X1_14 ( );
FILL FILL_1_AOI22X1_14 ( );
FILL FILL_2_AOI22X1_14 ( );
FILL FILL_3_AOI22X1_14 ( );
FILL FILL_4_AOI22X1_14 ( );
FILL FILL_5_AOI22X1_14 ( );
FILL FILL_6_AOI22X1_14 ( );
FILL FILL_7_AOI22X1_14 ( );
FILL FILL_8_AOI22X1_14 ( );
FILL FILL_9_AOI22X1_14 ( );
FILL FILL_10_AOI22X1_14 ( );
FILL FILL_11_AOI22X1_14 ( );
FILL FILL_0_INVX1_88 ( );
FILL FILL_1_INVX1_88 ( );
FILL FILL_2_INVX1_88 ( );
FILL FILL_3_INVX1_88 ( );
FILL FILL_4_INVX1_88 ( );
FILL FILL_0_DFFSR_235 ( );
FILL FILL_1_DFFSR_235 ( );
FILL FILL_2_DFFSR_235 ( );
FILL FILL_3_DFFSR_235 ( );
FILL FILL_4_DFFSR_235 ( );
FILL FILL_5_DFFSR_235 ( );
FILL FILL_6_DFFSR_235 ( );
FILL FILL_7_DFFSR_235 ( );
FILL FILL_8_DFFSR_235 ( );
FILL FILL_9_DFFSR_235 ( );
FILL FILL_10_DFFSR_235 ( );
FILL FILL_11_DFFSR_235 ( );
FILL FILL_12_DFFSR_235 ( );
FILL FILL_13_DFFSR_235 ( );
FILL FILL_14_DFFSR_235 ( );
FILL FILL_15_DFFSR_235 ( );
FILL FILL_16_DFFSR_235 ( );
FILL FILL_17_DFFSR_235 ( );
FILL FILL_18_DFFSR_235 ( );
FILL FILL_19_DFFSR_235 ( );
FILL FILL_20_DFFSR_235 ( );
FILL FILL_21_DFFSR_235 ( );
FILL FILL_22_DFFSR_235 ( );
FILL FILL_23_DFFSR_235 ( );
FILL FILL_24_DFFSR_235 ( );
FILL FILL_25_DFFSR_235 ( );
FILL FILL_26_DFFSR_235 ( );
FILL FILL_27_DFFSR_235 ( );
FILL FILL_28_DFFSR_235 ( );
FILL FILL_29_DFFSR_235 ( );
FILL FILL_30_DFFSR_235 ( );
FILL FILL_31_DFFSR_235 ( );
FILL FILL_32_DFFSR_235 ( );
FILL FILL_33_DFFSR_235 ( );
FILL FILL_34_DFFSR_235 ( );
FILL FILL_35_DFFSR_235 ( );
FILL FILL_36_DFFSR_235 ( );
FILL FILL_37_DFFSR_235 ( );
FILL FILL_38_DFFSR_235 ( );
FILL FILL_39_DFFSR_235 ( );
FILL FILL_40_DFFSR_235 ( );
FILL FILL_41_DFFSR_235 ( );
FILL FILL_42_DFFSR_235 ( );
FILL FILL_43_DFFSR_235 ( );
FILL FILL_44_DFFSR_235 ( );
FILL FILL_45_DFFSR_235 ( );
FILL FILL_46_DFFSR_235 ( );
FILL FILL_47_DFFSR_235 ( );
FILL FILL_48_DFFSR_235 ( );
FILL FILL_49_DFFSR_235 ( );
FILL FILL_50_DFFSR_235 ( );
FILL FILL_51_DFFSR_235 ( );
FILL FILL_0_BUFX2_67 ( );
FILL FILL_1_BUFX2_67 ( );
FILL FILL_2_BUFX2_67 ( );
FILL FILL_3_BUFX2_67 ( );
FILL FILL_4_BUFX2_67 ( );
FILL FILL_5_BUFX2_67 ( );
FILL FILL_6_BUFX2_67 ( );
FILL FILL_0_INVX1_66 ( );
FILL FILL_1_INVX1_66 ( );
FILL FILL_2_INVX1_66 ( );
FILL FILL_3_INVX1_66 ( );
FILL FILL_4_INVX1_66 ( );
FILL FILL_0_AOI22X1_9 ( );
FILL FILL_1_AOI22X1_9 ( );
FILL FILL_2_AOI22X1_9 ( );
FILL FILL_3_AOI22X1_9 ( );
FILL FILL_4_AOI22X1_9 ( );
FILL FILL_5_AOI22X1_9 ( );
FILL FILL_6_AOI22X1_9 ( );
FILL FILL_7_AOI22X1_9 ( );
FILL FILL_8_AOI22X1_9 ( );
FILL FILL_9_AOI22X1_9 ( );
FILL FILL_10_AOI22X1_9 ( );
FILL FILL_11_AOI22X1_9 ( );
FILL FILL_0_OAI22X1_27 ( );
FILL FILL_1_OAI22X1_27 ( );
FILL FILL_2_OAI22X1_27 ( );
FILL FILL_3_OAI22X1_27 ( );
FILL FILL_4_OAI22X1_27 ( );
FILL FILL_5_OAI22X1_27 ( );
FILL FILL_6_OAI22X1_27 ( );
FILL FILL_7_OAI22X1_27 ( );
FILL FILL_8_OAI22X1_27 ( );
FILL FILL_9_OAI22X1_27 ( );
FILL FILL_10_OAI22X1_27 ( );
FILL FILL_0_NOR2X1_35 ( );
FILL FILL_1_NOR2X1_35 ( );
FILL FILL_2_NOR2X1_35 ( );
FILL FILL_3_NOR2X1_35 ( );
FILL FILL_4_NOR2X1_35 ( );
FILL FILL_5_NOR2X1_35 ( );
FILL FILL_6_NOR2X1_35 ( );
FILL FILL_0_DFFSR_143 ( );
FILL FILL_1_DFFSR_143 ( );
FILL FILL_2_DFFSR_143 ( );
FILL FILL_3_DFFSR_143 ( );
FILL FILL_4_DFFSR_143 ( );
FILL FILL_5_DFFSR_143 ( );
FILL FILL_6_DFFSR_143 ( );
FILL FILL_7_DFFSR_143 ( );
FILL FILL_8_DFFSR_143 ( );
FILL FILL_9_DFFSR_143 ( );
FILL FILL_10_DFFSR_143 ( );
FILL FILL_11_DFFSR_143 ( );
FILL FILL_12_DFFSR_143 ( );
FILL FILL_13_DFFSR_143 ( );
FILL FILL_14_DFFSR_143 ( );
FILL FILL_15_DFFSR_143 ( );
FILL FILL_16_DFFSR_143 ( );
FILL FILL_17_DFFSR_143 ( );
FILL FILL_18_DFFSR_143 ( );
FILL FILL_19_DFFSR_143 ( );
FILL FILL_20_DFFSR_143 ( );
FILL FILL_21_DFFSR_143 ( );
FILL FILL_22_DFFSR_143 ( );
FILL FILL_23_DFFSR_143 ( );
FILL FILL_24_DFFSR_143 ( );
FILL FILL_25_DFFSR_143 ( );
FILL FILL_26_DFFSR_143 ( );
FILL FILL_27_DFFSR_143 ( );
FILL FILL_28_DFFSR_143 ( );
FILL FILL_29_DFFSR_143 ( );
FILL FILL_30_DFFSR_143 ( );
FILL FILL_31_DFFSR_143 ( );
FILL FILL_32_DFFSR_143 ( );
FILL FILL_33_DFFSR_143 ( );
FILL FILL_34_DFFSR_143 ( );
FILL FILL_35_DFFSR_143 ( );
FILL FILL_36_DFFSR_143 ( );
FILL FILL_37_DFFSR_143 ( );
FILL FILL_38_DFFSR_143 ( );
FILL FILL_39_DFFSR_143 ( );
FILL FILL_40_DFFSR_143 ( );
FILL FILL_41_DFFSR_143 ( );
FILL FILL_42_DFFSR_143 ( );
FILL FILL_43_DFFSR_143 ( );
FILL FILL_44_DFFSR_143 ( );
FILL FILL_45_DFFSR_143 ( );
FILL FILL_46_DFFSR_143 ( );
FILL FILL_47_DFFSR_143 ( );
FILL FILL_48_DFFSR_143 ( );
FILL FILL_49_DFFSR_143 ( );
FILL FILL_50_DFFSR_143 ( );
FILL FILL_51_DFFSR_143 ( );
FILL FILL_0_DFFSR_167 ( );
FILL FILL_1_DFFSR_167 ( );
FILL FILL_2_DFFSR_167 ( );
FILL FILL_3_DFFSR_167 ( );
FILL FILL_4_DFFSR_167 ( );
FILL FILL_5_DFFSR_167 ( );
FILL FILL_6_DFFSR_167 ( );
FILL FILL_7_DFFSR_167 ( );
FILL FILL_8_DFFSR_167 ( );
FILL FILL_9_DFFSR_167 ( );
FILL FILL_10_DFFSR_167 ( );
FILL FILL_11_DFFSR_167 ( );
FILL FILL_12_DFFSR_167 ( );
FILL FILL_13_DFFSR_167 ( );
FILL FILL_14_DFFSR_167 ( );
FILL FILL_15_DFFSR_167 ( );
FILL FILL_16_DFFSR_167 ( );
FILL FILL_17_DFFSR_167 ( );
FILL FILL_18_DFFSR_167 ( );
FILL FILL_19_DFFSR_167 ( );
FILL FILL_20_DFFSR_167 ( );
FILL FILL_21_DFFSR_167 ( );
FILL FILL_22_DFFSR_167 ( );
FILL FILL_23_DFFSR_167 ( );
FILL FILL_24_DFFSR_167 ( );
FILL FILL_25_DFFSR_167 ( );
FILL FILL_26_DFFSR_167 ( );
FILL FILL_27_DFFSR_167 ( );
FILL FILL_28_DFFSR_167 ( );
FILL FILL_29_DFFSR_167 ( );
FILL FILL_30_DFFSR_167 ( );
FILL FILL_31_DFFSR_167 ( );
FILL FILL_32_DFFSR_167 ( );
FILL FILL_33_DFFSR_167 ( );
FILL FILL_34_DFFSR_167 ( );
FILL FILL_35_DFFSR_167 ( );
FILL FILL_36_DFFSR_167 ( );
FILL FILL_37_DFFSR_167 ( );
FILL FILL_38_DFFSR_167 ( );
FILL FILL_39_DFFSR_167 ( );
FILL FILL_40_DFFSR_167 ( );
FILL FILL_41_DFFSR_167 ( );
FILL FILL_42_DFFSR_167 ( );
FILL FILL_43_DFFSR_167 ( );
FILL FILL_44_DFFSR_167 ( );
FILL FILL_45_DFFSR_167 ( );
FILL FILL_46_DFFSR_167 ( );
FILL FILL_47_DFFSR_167 ( );
FILL FILL_48_DFFSR_167 ( );
FILL FILL_49_DFFSR_167 ( );
FILL FILL_50_DFFSR_167 ( );
FILL FILL_51_DFFSR_167 ( );
FILL FILL_0_INVX1_157 ( );
FILL FILL_1_INVX1_157 ( );
FILL FILL_2_INVX1_157 ( );
FILL FILL_3_INVX1_157 ( );
FILL FILL_4_INVX1_157 ( );
FILL FILL_0_NAND3X1_185 ( );
FILL FILL_1_NAND3X1_185 ( );
FILL FILL_2_NAND3X1_185 ( );
FILL FILL_3_NAND3X1_185 ( );
FILL FILL_4_NAND3X1_185 ( );
FILL FILL_5_NAND3X1_185 ( );
FILL FILL_6_NAND3X1_185 ( );
FILL FILL_7_NAND3X1_185 ( );
FILL FILL_8_NAND3X1_185 ( );
FILL FILL_0_NAND3X1_187 ( );
FILL FILL_1_NAND3X1_187 ( );
FILL FILL_2_NAND3X1_187 ( );
FILL FILL_3_NAND3X1_187 ( );
FILL FILL_4_NAND3X1_187 ( );
FILL FILL_5_NAND3X1_187 ( );
FILL FILL_6_NAND3X1_187 ( );
FILL FILL_7_NAND3X1_187 ( );
FILL FILL_8_NAND3X1_187 ( );
FILL FILL_0_INVX1_204 ( );
FILL FILL_1_INVX1_204 ( );
FILL FILL_2_INVX1_204 ( );
FILL FILL_3_INVX1_204 ( );
FILL FILL_4_INVX1_204 ( );
FILL FILL_0_NAND3X1_137 ( );
FILL FILL_1_NAND3X1_137 ( );
FILL FILL_2_NAND3X1_137 ( );
FILL FILL_3_NAND3X1_137 ( );
FILL FILL_4_NAND3X1_137 ( );
FILL FILL_5_NAND3X1_137 ( );
FILL FILL_6_NAND3X1_137 ( );
FILL FILL_7_NAND3X1_137 ( );
FILL FILL_8_NAND3X1_137 ( );
FILL FILL_9_NAND3X1_137 ( );
FILL FILL_0_NOR3X1_5 ( );
FILL FILL_1_NOR3X1_5 ( );
FILL FILL_2_NOR3X1_5 ( );
FILL FILL_3_NOR3X1_5 ( );
FILL FILL_4_NOR3X1_5 ( );
FILL FILL_5_NOR3X1_5 ( );
FILL FILL_6_NOR3X1_5 ( );
FILL FILL_7_NOR3X1_5 ( );
FILL FILL_8_NOR3X1_5 ( );
FILL FILL_9_NOR3X1_5 ( );
FILL FILL_10_NOR3X1_5 ( );
FILL FILL_11_NOR3X1_5 ( );
FILL FILL_12_NOR3X1_5 ( );
FILL FILL_13_NOR3X1_5 ( );
FILL FILL_14_NOR3X1_5 ( );
FILL FILL_15_NOR3X1_5 ( );
FILL FILL_16_NOR3X1_5 ( );
FILL FILL_17_NOR3X1_5 ( );
FILL FILL_18_NOR3X1_5 ( );
FILL FILL_0_NAND3X1_154 ( );
FILL FILL_1_NAND3X1_154 ( );
FILL FILL_2_NAND3X1_154 ( );
FILL FILL_3_NAND3X1_154 ( );
FILL FILL_4_NAND3X1_154 ( );
FILL FILL_5_NAND3X1_154 ( );
FILL FILL_6_NAND3X1_154 ( );
FILL FILL_7_NAND3X1_154 ( );
FILL FILL_8_NAND3X1_154 ( );
FILL FILL_9_NAND3X1_154 ( );
FILL FILL_0_INVX1_148 ( );
FILL FILL_1_INVX1_148 ( );
FILL FILL_2_INVX1_148 ( );
FILL FILL_3_INVX1_148 ( );
FILL FILL_0_INVX1_147 ( );
FILL FILL_1_INVX1_147 ( );
FILL FILL_2_INVX1_147 ( );
FILL FILL_3_INVX1_147 ( );
FILL FILL_4_INVX1_147 ( );
FILL FILL_0_NAND3X1_155 ( );
FILL FILL_1_NAND3X1_155 ( );
FILL FILL_2_NAND3X1_155 ( );
FILL FILL_3_NAND3X1_155 ( );
FILL FILL_4_NAND3X1_155 ( );
FILL FILL_5_NAND3X1_155 ( );
FILL FILL_6_NAND3X1_155 ( );
FILL FILL_7_NAND3X1_155 ( );
FILL FILL_8_NAND3X1_155 ( );
FILL FILL_0_OAI21X1_35 ( );
FILL FILL_1_OAI21X1_35 ( );
FILL FILL_2_OAI21X1_35 ( );
FILL FILL_3_OAI21X1_35 ( );
FILL FILL_4_OAI21X1_35 ( );
FILL FILL_5_OAI21X1_35 ( );
FILL FILL_6_OAI21X1_35 ( );
FILL FILL_7_OAI21X1_35 ( );
FILL FILL_8_OAI21X1_35 ( );
FILL FILL_0_BUFX2_53 ( );
FILL FILL_1_BUFX2_53 ( );
FILL FILL_2_BUFX2_53 ( );
FILL FILL_3_BUFX2_53 ( );
FILL FILL_4_BUFX2_53 ( );
FILL FILL_5_BUFX2_53 ( );
FILL FILL_6_BUFX2_53 ( );
FILL FILL_0_OAI21X1_95 ( );
FILL FILL_1_OAI21X1_95 ( );
FILL FILL_2_OAI21X1_95 ( );
FILL FILL_3_OAI21X1_95 ( );
FILL FILL_4_OAI21X1_95 ( );
FILL FILL_5_OAI21X1_95 ( );
FILL FILL_6_OAI21X1_95 ( );
FILL FILL_7_OAI21X1_95 ( );
FILL FILL_8_OAI21X1_95 ( );
FILL FILL_9_OAI21X1_95 ( );
FILL FILL_0_INVX1_131 ( );
FILL FILL_1_INVX1_131 ( );
FILL FILL_2_INVX1_131 ( );
FILL FILL_3_INVX1_131 ( );
FILL FILL_0_NAND2X1_170 ( );
FILL FILL_1_NAND2X1_170 ( );
FILL FILL_2_NAND2X1_170 ( );
FILL FILL_3_NAND2X1_170 ( );
FILL FILL_4_NAND2X1_170 ( );
FILL FILL_5_NAND2X1_170 ( );
FILL FILL_6_NAND2X1_170 ( );
FILL FILL_0_AOI21X1_49 ( );
FILL FILL_1_AOI21X1_49 ( );
FILL FILL_2_AOI21X1_49 ( );
FILL FILL_3_AOI21X1_49 ( );
FILL FILL_4_AOI21X1_49 ( );
FILL FILL_5_AOI21X1_49 ( );
FILL FILL_6_AOI21X1_49 ( );
FILL FILL_7_AOI21X1_49 ( );
FILL FILL_8_AOI21X1_49 ( );
FILL FILL_0_DFFSR_204 ( );
FILL FILL_1_DFFSR_204 ( );
FILL FILL_2_DFFSR_204 ( );
FILL FILL_3_DFFSR_204 ( );
FILL FILL_4_DFFSR_204 ( );
FILL FILL_5_DFFSR_204 ( );
FILL FILL_6_DFFSR_204 ( );
FILL FILL_7_DFFSR_204 ( );
FILL FILL_8_DFFSR_204 ( );
FILL FILL_9_DFFSR_204 ( );
FILL FILL_10_DFFSR_204 ( );
FILL FILL_11_DFFSR_204 ( );
FILL FILL_12_DFFSR_204 ( );
FILL FILL_13_DFFSR_204 ( );
FILL FILL_14_DFFSR_204 ( );
FILL FILL_15_DFFSR_204 ( );
FILL FILL_16_DFFSR_204 ( );
FILL FILL_17_DFFSR_204 ( );
FILL FILL_18_DFFSR_204 ( );
FILL FILL_19_DFFSR_204 ( );
FILL FILL_20_DFFSR_204 ( );
FILL FILL_21_DFFSR_204 ( );
FILL FILL_22_DFFSR_204 ( );
FILL FILL_23_DFFSR_204 ( );
FILL FILL_24_DFFSR_204 ( );
FILL FILL_25_DFFSR_204 ( );
FILL FILL_26_DFFSR_204 ( );
FILL FILL_27_DFFSR_204 ( );
FILL FILL_28_DFFSR_204 ( );
FILL FILL_29_DFFSR_204 ( );
FILL FILL_30_DFFSR_204 ( );
FILL FILL_31_DFFSR_204 ( );
FILL FILL_32_DFFSR_204 ( );
FILL FILL_33_DFFSR_204 ( );
FILL FILL_34_DFFSR_204 ( );
FILL FILL_35_DFFSR_204 ( );
FILL FILL_36_DFFSR_204 ( );
FILL FILL_37_DFFSR_204 ( );
FILL FILL_38_DFFSR_204 ( );
FILL FILL_39_DFFSR_204 ( );
FILL FILL_40_DFFSR_204 ( );
FILL FILL_41_DFFSR_204 ( );
FILL FILL_42_DFFSR_204 ( );
FILL FILL_43_DFFSR_204 ( );
FILL FILL_44_DFFSR_204 ( );
FILL FILL_45_DFFSR_204 ( );
FILL FILL_46_DFFSR_204 ( );
FILL FILL_47_DFFSR_204 ( );
FILL FILL_48_DFFSR_204 ( );
FILL FILL_49_DFFSR_204 ( );
FILL FILL_50_DFFSR_204 ( );
FILL FILL_0_DFFSR_198 ( );
FILL FILL_1_DFFSR_198 ( );
FILL FILL_2_DFFSR_198 ( );
FILL FILL_3_DFFSR_198 ( );
FILL FILL_4_DFFSR_198 ( );
FILL FILL_5_DFFSR_198 ( );
FILL FILL_6_DFFSR_198 ( );
FILL FILL_7_DFFSR_198 ( );
FILL FILL_8_DFFSR_198 ( );
FILL FILL_9_DFFSR_198 ( );
FILL FILL_10_DFFSR_198 ( );
FILL FILL_11_DFFSR_198 ( );
FILL FILL_12_DFFSR_198 ( );
FILL FILL_13_DFFSR_198 ( );
FILL FILL_14_DFFSR_198 ( );
FILL FILL_15_DFFSR_198 ( );
FILL FILL_16_DFFSR_198 ( );
FILL FILL_17_DFFSR_198 ( );
FILL FILL_18_DFFSR_198 ( );
FILL FILL_19_DFFSR_198 ( );
FILL FILL_20_DFFSR_198 ( );
FILL FILL_21_DFFSR_198 ( );
FILL FILL_22_DFFSR_198 ( );
FILL FILL_23_DFFSR_198 ( );
FILL FILL_24_DFFSR_198 ( );
FILL FILL_25_DFFSR_198 ( );
FILL FILL_26_DFFSR_198 ( );
FILL FILL_27_DFFSR_198 ( );
FILL FILL_28_DFFSR_198 ( );
FILL FILL_29_DFFSR_198 ( );
FILL FILL_30_DFFSR_198 ( );
FILL FILL_31_DFFSR_198 ( );
FILL FILL_32_DFFSR_198 ( );
FILL FILL_33_DFFSR_198 ( );
FILL FILL_34_DFFSR_198 ( );
FILL FILL_35_DFFSR_198 ( );
FILL FILL_36_DFFSR_198 ( );
FILL FILL_37_DFFSR_198 ( );
FILL FILL_38_DFFSR_198 ( );
FILL FILL_39_DFFSR_198 ( );
FILL FILL_40_DFFSR_198 ( );
FILL FILL_41_DFFSR_198 ( );
FILL FILL_42_DFFSR_198 ( );
FILL FILL_43_DFFSR_198 ( );
FILL FILL_44_DFFSR_198 ( );
FILL FILL_45_DFFSR_198 ( );
FILL FILL_46_DFFSR_198 ( );
FILL FILL_47_DFFSR_198 ( );
FILL FILL_48_DFFSR_198 ( );
FILL FILL_49_DFFSR_198 ( );
FILL FILL_50_DFFSR_198 ( );
FILL FILL_0_DFFSR_211 ( );
FILL FILL_1_DFFSR_211 ( );
FILL FILL_2_DFFSR_211 ( );
FILL FILL_3_DFFSR_211 ( );
FILL FILL_4_DFFSR_211 ( );
FILL FILL_5_DFFSR_211 ( );
FILL FILL_6_DFFSR_211 ( );
FILL FILL_7_DFFSR_211 ( );
FILL FILL_8_DFFSR_211 ( );
FILL FILL_9_DFFSR_211 ( );
FILL FILL_10_DFFSR_211 ( );
FILL FILL_11_DFFSR_211 ( );
FILL FILL_12_DFFSR_211 ( );
FILL FILL_13_DFFSR_211 ( );
FILL FILL_14_DFFSR_211 ( );
FILL FILL_15_DFFSR_211 ( );
FILL FILL_16_DFFSR_211 ( );
FILL FILL_17_DFFSR_211 ( );
FILL FILL_18_DFFSR_211 ( );
FILL FILL_19_DFFSR_211 ( );
FILL FILL_20_DFFSR_211 ( );
FILL FILL_21_DFFSR_211 ( );
FILL FILL_22_DFFSR_211 ( );
FILL FILL_23_DFFSR_211 ( );
FILL FILL_24_DFFSR_211 ( );
FILL FILL_25_DFFSR_211 ( );
FILL FILL_26_DFFSR_211 ( );
FILL FILL_27_DFFSR_211 ( );
FILL FILL_28_DFFSR_211 ( );
FILL FILL_29_DFFSR_211 ( );
FILL FILL_30_DFFSR_211 ( );
FILL FILL_31_DFFSR_211 ( );
FILL FILL_32_DFFSR_211 ( );
FILL FILL_33_DFFSR_211 ( );
FILL FILL_34_DFFSR_211 ( );
FILL FILL_35_DFFSR_211 ( );
FILL FILL_36_DFFSR_211 ( );
FILL FILL_37_DFFSR_211 ( );
FILL FILL_38_DFFSR_211 ( );
FILL FILL_39_DFFSR_211 ( );
FILL FILL_40_DFFSR_211 ( );
FILL FILL_41_DFFSR_211 ( );
FILL FILL_42_DFFSR_211 ( );
FILL FILL_43_DFFSR_211 ( );
FILL FILL_44_DFFSR_211 ( );
FILL FILL_45_DFFSR_211 ( );
FILL FILL_46_DFFSR_211 ( );
FILL FILL_47_DFFSR_211 ( );
FILL FILL_48_DFFSR_211 ( );
FILL FILL_49_DFFSR_211 ( );
FILL FILL_50_DFFSR_211 ( );
FILL FILL_51_DFFSR_211 ( );
FILL FILL_0_NOR3X1_3 ( );
FILL FILL_1_NOR3X1_3 ( );
FILL FILL_2_NOR3X1_3 ( );
FILL FILL_3_NOR3X1_3 ( );
FILL FILL_4_NOR3X1_3 ( );
FILL FILL_5_NOR3X1_3 ( );
FILL FILL_6_NOR3X1_3 ( );
FILL FILL_7_NOR3X1_3 ( );
FILL FILL_8_NOR3X1_3 ( );
FILL FILL_9_NOR3X1_3 ( );
FILL FILL_10_NOR3X1_3 ( );
FILL FILL_11_NOR3X1_3 ( );
FILL FILL_12_NOR3X1_3 ( );
FILL FILL_13_NOR3X1_3 ( );
FILL FILL_14_NOR3X1_3 ( );
FILL FILL_15_NOR3X1_3 ( );
FILL FILL_16_NOR3X1_3 ( );
FILL FILL_17_NOR3X1_3 ( );
FILL FILL_0_OAI22X1_36 ( );
FILL FILL_1_OAI22X1_36 ( );
FILL FILL_2_OAI22X1_36 ( );
FILL FILL_3_OAI22X1_36 ( );
FILL FILL_4_OAI22X1_36 ( );
FILL FILL_5_OAI22X1_36 ( );
FILL FILL_6_OAI22X1_36 ( );
FILL FILL_7_OAI22X1_36 ( );
FILL FILL_8_OAI22X1_36 ( );
FILL FILL_9_OAI22X1_36 ( );
FILL FILL_10_OAI22X1_36 ( );
FILL FILL_11_OAI22X1_36 ( );
FILL FILL_0_NAND2X1_37 ( );
FILL FILL_1_NAND2X1_37 ( );
FILL FILL_2_NAND2X1_37 ( );
FILL FILL_3_NAND2X1_37 ( );
FILL FILL_4_NAND2X1_37 ( );
FILL FILL_5_NAND2X1_37 ( );
FILL FILL_6_NAND2X1_37 ( );
FILL FILL_0_NAND3X1_68 ( );
FILL FILL_1_NAND3X1_68 ( );
FILL FILL_2_NAND3X1_68 ( );
FILL FILL_3_NAND3X1_68 ( );
FILL FILL_4_NAND3X1_68 ( );
FILL FILL_5_NAND3X1_68 ( );
FILL FILL_6_NAND3X1_68 ( );
FILL FILL_7_NAND3X1_68 ( );
FILL FILL_8_NAND3X1_68 ( );
FILL FILL_0_AND2X2_19 ( );
FILL FILL_1_AND2X2_19 ( );
FILL FILL_2_AND2X2_19 ( );
FILL FILL_3_AND2X2_19 ( );
FILL FILL_4_AND2X2_19 ( );
FILL FILL_5_AND2X2_19 ( );
FILL FILL_6_AND2X2_19 ( );
FILL FILL_7_AND2X2_19 ( );
FILL FILL_8_AND2X2_19 ( );
FILL FILL_9_AND2X2_19 ( );
FILL FILL_0_NOR2X1_37 ( );
FILL FILL_1_NOR2X1_37 ( );
FILL FILL_2_NOR2X1_37 ( );
FILL FILL_3_NOR2X1_37 ( );
FILL FILL_4_NOR2X1_37 ( );
FILL FILL_5_NOR2X1_37 ( );
FILL FILL_6_NOR2X1_37 ( );
FILL FILL_0_NAND3X1_71 ( );
FILL FILL_1_NAND3X1_71 ( );
FILL FILL_2_NAND3X1_71 ( );
FILL FILL_3_NAND3X1_71 ( );
FILL FILL_4_NAND3X1_71 ( );
FILL FILL_5_NAND3X1_71 ( );
FILL FILL_6_NAND3X1_71 ( );
FILL FILL_7_NAND3X1_71 ( );
FILL FILL_8_NAND3X1_71 ( );
FILL FILL_0_NAND3X1_69 ( );
FILL FILL_1_NAND3X1_69 ( );
FILL FILL_2_NAND3X1_69 ( );
FILL FILL_3_NAND3X1_69 ( );
FILL FILL_4_NAND3X1_69 ( );
FILL FILL_5_NAND3X1_69 ( );
FILL FILL_6_NAND3X1_69 ( );
FILL FILL_7_NAND3X1_69 ( );
FILL FILL_8_NAND3X1_69 ( );
FILL FILL_0_DFFSR_137 ( );
FILL FILL_1_DFFSR_137 ( );
FILL FILL_2_DFFSR_137 ( );
FILL FILL_3_DFFSR_137 ( );
FILL FILL_4_DFFSR_137 ( );
FILL FILL_5_DFFSR_137 ( );
FILL FILL_6_DFFSR_137 ( );
FILL FILL_7_DFFSR_137 ( );
FILL FILL_8_DFFSR_137 ( );
FILL FILL_9_DFFSR_137 ( );
FILL FILL_10_DFFSR_137 ( );
FILL FILL_11_DFFSR_137 ( );
FILL FILL_12_DFFSR_137 ( );
FILL FILL_13_DFFSR_137 ( );
FILL FILL_14_DFFSR_137 ( );
FILL FILL_15_DFFSR_137 ( );
FILL FILL_16_DFFSR_137 ( );
FILL FILL_17_DFFSR_137 ( );
FILL FILL_18_DFFSR_137 ( );
FILL FILL_19_DFFSR_137 ( );
FILL FILL_20_DFFSR_137 ( );
FILL FILL_21_DFFSR_137 ( );
FILL FILL_22_DFFSR_137 ( );
FILL FILL_23_DFFSR_137 ( );
FILL FILL_24_DFFSR_137 ( );
FILL FILL_25_DFFSR_137 ( );
FILL FILL_26_DFFSR_137 ( );
FILL FILL_27_DFFSR_137 ( );
FILL FILL_28_DFFSR_137 ( );
FILL FILL_29_DFFSR_137 ( );
FILL FILL_30_DFFSR_137 ( );
FILL FILL_31_DFFSR_137 ( );
FILL FILL_32_DFFSR_137 ( );
FILL FILL_33_DFFSR_137 ( );
FILL FILL_34_DFFSR_137 ( );
FILL FILL_35_DFFSR_137 ( );
FILL FILL_36_DFFSR_137 ( );
FILL FILL_37_DFFSR_137 ( );
FILL FILL_38_DFFSR_137 ( );
FILL FILL_39_DFFSR_137 ( );
FILL FILL_40_DFFSR_137 ( );
FILL FILL_41_DFFSR_137 ( );
FILL FILL_42_DFFSR_137 ( );
FILL FILL_43_DFFSR_137 ( );
FILL FILL_44_DFFSR_137 ( );
FILL FILL_45_DFFSR_137 ( );
FILL FILL_46_DFFSR_137 ( );
FILL FILL_47_DFFSR_137 ( );
FILL FILL_48_DFFSR_137 ( );
FILL FILL_49_DFFSR_137 ( );
FILL FILL_50_DFFSR_137 ( );
FILL FILL_51_DFFSR_137 ( );
FILL FILL_0_INVX1_95 ( );
FILL FILL_1_INVX1_95 ( );
FILL FILL_2_INVX1_95 ( );
FILL FILL_3_INVX1_95 ( );
FILL FILL_4_INVX1_95 ( );
FILL FILL_0_DFFSR_216 ( );
FILL FILL_1_DFFSR_216 ( );
FILL FILL_2_DFFSR_216 ( );
FILL FILL_3_DFFSR_216 ( );
FILL FILL_4_DFFSR_216 ( );
FILL FILL_5_DFFSR_216 ( );
FILL FILL_6_DFFSR_216 ( );
FILL FILL_7_DFFSR_216 ( );
FILL FILL_8_DFFSR_216 ( );
FILL FILL_9_DFFSR_216 ( );
FILL FILL_10_DFFSR_216 ( );
FILL FILL_11_DFFSR_216 ( );
FILL FILL_12_DFFSR_216 ( );
FILL FILL_13_DFFSR_216 ( );
FILL FILL_14_DFFSR_216 ( );
FILL FILL_15_DFFSR_216 ( );
FILL FILL_16_DFFSR_216 ( );
FILL FILL_17_DFFSR_216 ( );
FILL FILL_18_DFFSR_216 ( );
FILL FILL_19_DFFSR_216 ( );
FILL FILL_20_DFFSR_216 ( );
FILL FILL_21_DFFSR_216 ( );
FILL FILL_22_DFFSR_216 ( );
FILL FILL_23_DFFSR_216 ( );
FILL FILL_24_DFFSR_216 ( );
FILL FILL_25_DFFSR_216 ( );
FILL FILL_26_DFFSR_216 ( );
FILL FILL_27_DFFSR_216 ( );
FILL FILL_28_DFFSR_216 ( );
FILL FILL_29_DFFSR_216 ( );
FILL FILL_30_DFFSR_216 ( );
FILL FILL_31_DFFSR_216 ( );
FILL FILL_32_DFFSR_216 ( );
FILL FILL_33_DFFSR_216 ( );
FILL FILL_34_DFFSR_216 ( );
FILL FILL_35_DFFSR_216 ( );
FILL FILL_36_DFFSR_216 ( );
FILL FILL_37_DFFSR_216 ( );
FILL FILL_38_DFFSR_216 ( );
FILL FILL_39_DFFSR_216 ( );
FILL FILL_40_DFFSR_216 ( );
FILL FILL_41_DFFSR_216 ( );
FILL FILL_42_DFFSR_216 ( );
FILL FILL_43_DFFSR_216 ( );
FILL FILL_44_DFFSR_216 ( );
FILL FILL_45_DFFSR_216 ( );
FILL FILL_46_DFFSR_216 ( );
FILL FILL_47_DFFSR_216 ( );
FILL FILL_48_DFFSR_216 ( );
FILL FILL_49_DFFSR_216 ( );
FILL FILL_50_DFFSR_216 ( );
FILL FILL_0_NAND3X1_186 ( );
FILL FILL_1_NAND3X1_186 ( );
FILL FILL_2_NAND3X1_186 ( );
FILL FILL_3_NAND3X1_186 ( );
FILL FILL_4_NAND3X1_186 ( );
FILL FILL_5_NAND3X1_186 ( );
FILL FILL_6_NAND3X1_186 ( );
FILL FILL_7_NAND3X1_186 ( );
FILL FILL_8_NAND3X1_186 ( );
FILL FILL_0_NAND3X1_189 ( );
FILL FILL_1_NAND3X1_189 ( );
FILL FILL_2_NAND3X1_189 ( );
FILL FILL_3_NAND3X1_189 ( );
FILL FILL_4_NAND3X1_189 ( );
FILL FILL_5_NAND3X1_189 ( );
FILL FILL_6_NAND3X1_189 ( );
FILL FILL_7_NAND3X1_189 ( );
FILL FILL_8_NAND3X1_189 ( );
FILL FILL_0_NAND3X1_188 ( );
FILL FILL_1_NAND3X1_188 ( );
FILL FILL_2_NAND3X1_188 ( );
FILL FILL_3_NAND3X1_188 ( );
FILL FILL_4_NAND3X1_188 ( );
FILL FILL_5_NAND3X1_188 ( );
FILL FILL_6_NAND3X1_188 ( );
FILL FILL_7_NAND3X1_188 ( );
FILL FILL_8_NAND3X1_188 ( );
FILL FILL_9_NAND3X1_188 ( );
FILL FILL_0_NAND3X1_190 ( );
FILL FILL_1_NAND3X1_190 ( );
FILL FILL_2_NAND3X1_190 ( );
FILL FILL_3_NAND3X1_190 ( );
FILL FILL_4_NAND3X1_190 ( );
FILL FILL_5_NAND3X1_190 ( );
FILL FILL_6_NAND3X1_190 ( );
FILL FILL_7_NAND3X1_190 ( );
FILL FILL_8_NAND3X1_190 ( );
FILL FILL_0_NAND3X1_191 ( );
FILL FILL_1_NAND3X1_191 ( );
FILL FILL_2_NAND3X1_191 ( );
FILL FILL_3_NAND3X1_191 ( );
FILL FILL_4_NAND3X1_191 ( );
FILL FILL_5_NAND3X1_191 ( );
FILL FILL_6_NAND3X1_191 ( );
FILL FILL_7_NAND3X1_191 ( );
FILL FILL_8_NAND3X1_191 ( );
FILL FILL_9_NAND3X1_191 ( );
FILL FILL_0_OAI21X1_42 ( );
FILL FILL_1_OAI21X1_42 ( );
FILL FILL_2_OAI21X1_42 ( );
FILL FILL_3_OAI21X1_42 ( );
FILL FILL_4_OAI21X1_42 ( );
FILL FILL_5_OAI21X1_42 ( );
FILL FILL_6_OAI21X1_42 ( );
FILL FILL_7_OAI21X1_42 ( );
FILL FILL_8_OAI21X1_42 ( );
FILL FILL_9_OAI21X1_42 ( );
FILL FILL_0_INVX1_149 ( );
FILL FILL_1_INVX1_149 ( );
FILL FILL_2_INVX1_149 ( );
FILL FILL_3_INVX1_149 ( );
FILL FILL_4_INVX1_149 ( );
FILL FILL_0_OAI21X1_34 ( );
FILL FILL_1_OAI21X1_34 ( );
FILL FILL_2_OAI21X1_34 ( );
FILL FILL_3_OAI21X1_34 ( );
FILL FILL_4_OAI21X1_34 ( );
FILL FILL_5_OAI21X1_34 ( );
FILL FILL_6_OAI21X1_34 ( );
FILL FILL_7_OAI21X1_34 ( );
FILL FILL_8_OAI21X1_34 ( );
FILL FILL_0_AOI21X1_17 ( );
FILL FILL_1_AOI21X1_17 ( );
FILL FILL_2_AOI21X1_17 ( );
FILL FILL_3_AOI21X1_17 ( );
FILL FILL_4_AOI21X1_17 ( );
FILL FILL_5_AOI21X1_17 ( );
FILL FILL_6_AOI21X1_17 ( );
FILL FILL_7_AOI21X1_17 ( );
FILL FILL_8_AOI21X1_17 ( );
FILL FILL_9_AOI21X1_17 ( );
FILL FILL_0_OAI21X1_43 ( );
FILL FILL_1_OAI21X1_43 ( );
FILL FILL_2_OAI21X1_43 ( );
FILL FILL_3_OAI21X1_43 ( );
FILL FILL_4_OAI21X1_43 ( );
FILL FILL_5_OAI21X1_43 ( );
FILL FILL_6_OAI21X1_43 ( );
FILL FILL_7_OAI21X1_43 ( );
FILL FILL_8_OAI21X1_43 ( );
FILL FILL_0_BUFX2_54 ( );
FILL FILL_1_BUFX2_54 ( );
FILL FILL_2_BUFX2_54 ( );
FILL FILL_3_BUFX2_54 ( );
FILL FILL_4_BUFX2_54 ( );
FILL FILL_5_BUFX2_54 ( );
FILL FILL_6_BUFX2_54 ( );
FILL FILL_0_BUFX2_39 ( );
FILL FILL_1_BUFX2_39 ( );
FILL FILL_2_BUFX2_39 ( );
FILL FILL_3_BUFX2_39 ( );
FILL FILL_4_BUFX2_39 ( );
FILL FILL_5_BUFX2_39 ( );
FILL FILL_6_BUFX2_39 ( );
FILL FILL_0_DFFPOSX1_39 ( );
FILL FILL_1_DFFPOSX1_39 ( );
FILL FILL_2_DFFPOSX1_39 ( );
FILL FILL_3_DFFPOSX1_39 ( );
FILL FILL_4_DFFPOSX1_39 ( );
FILL FILL_5_DFFPOSX1_39 ( );
FILL FILL_6_DFFPOSX1_39 ( );
FILL FILL_7_DFFPOSX1_39 ( );
FILL FILL_8_DFFPOSX1_39 ( );
FILL FILL_9_DFFPOSX1_39 ( );
FILL FILL_10_DFFPOSX1_39 ( );
FILL FILL_11_DFFPOSX1_39 ( );
FILL FILL_12_DFFPOSX1_39 ( );
FILL FILL_13_DFFPOSX1_39 ( );
FILL FILL_14_DFFPOSX1_39 ( );
FILL FILL_15_DFFPOSX1_39 ( );
FILL FILL_16_DFFPOSX1_39 ( );
FILL FILL_17_DFFPOSX1_39 ( );
FILL FILL_18_DFFPOSX1_39 ( );
FILL FILL_19_DFFPOSX1_39 ( );
FILL FILL_20_DFFPOSX1_39 ( );
FILL FILL_21_DFFPOSX1_39 ( );
FILL FILL_22_DFFPOSX1_39 ( );
FILL FILL_23_DFFPOSX1_39 ( );
FILL FILL_24_DFFPOSX1_39 ( );
FILL FILL_25_DFFPOSX1_39 ( );
FILL FILL_26_DFFPOSX1_39 ( );
FILL FILL_27_DFFPOSX1_39 ( );
FILL FILL_0_NAND2X1_146 ( );
FILL FILL_1_NAND2X1_146 ( );
FILL FILL_2_NAND2X1_146 ( );
FILL FILL_3_NAND2X1_146 ( );
FILL FILL_4_NAND2X1_146 ( );
FILL FILL_5_NAND2X1_146 ( );
FILL FILL_6_NAND2X1_146 ( );
FILL FILL_0_BUFX2_7 ( );
FILL FILL_1_BUFX2_7 ( );
FILL FILL_2_BUFX2_7 ( );
FILL FILL_3_BUFX2_7 ( );
FILL FILL_4_BUFX2_7 ( );
FILL FILL_5_BUFX2_7 ( );
FILL FILL_6_BUFX2_7 ( );
FILL FILL_0_NAND2X1_140 ( );
FILL FILL_1_NAND2X1_140 ( );
FILL FILL_2_NAND2X1_140 ( );
FILL FILL_3_NAND2X1_140 ( );
FILL FILL_4_NAND2X1_140 ( );
FILL FILL_5_NAND2X1_140 ( );
FILL FILL_6_NAND2X1_140 ( );
FILL FILL_0_AOI21X1_46 ( );
FILL FILL_1_AOI21X1_46 ( );
FILL FILL_2_AOI21X1_46 ( );
FILL FILL_3_AOI21X1_46 ( );
FILL FILL_4_AOI21X1_46 ( );
FILL FILL_5_AOI21X1_46 ( );
FILL FILL_6_AOI21X1_46 ( );
FILL FILL_7_AOI21X1_46 ( );
FILL FILL_8_AOI21X1_46 ( );
FILL FILL_0_DFFSR_220 ( );
FILL FILL_1_DFFSR_220 ( );
FILL FILL_2_DFFSR_220 ( );
FILL FILL_3_DFFSR_220 ( );
FILL FILL_4_DFFSR_220 ( );
FILL FILL_5_DFFSR_220 ( );
FILL FILL_6_DFFSR_220 ( );
FILL FILL_7_DFFSR_220 ( );
FILL FILL_8_DFFSR_220 ( );
FILL FILL_9_DFFSR_220 ( );
FILL FILL_10_DFFSR_220 ( );
FILL FILL_11_DFFSR_220 ( );
FILL FILL_12_DFFSR_220 ( );
FILL FILL_13_DFFSR_220 ( );
FILL FILL_14_DFFSR_220 ( );
FILL FILL_15_DFFSR_220 ( );
FILL FILL_16_DFFSR_220 ( );
FILL FILL_17_DFFSR_220 ( );
FILL FILL_18_DFFSR_220 ( );
FILL FILL_19_DFFSR_220 ( );
FILL FILL_20_DFFSR_220 ( );
FILL FILL_21_DFFSR_220 ( );
FILL FILL_22_DFFSR_220 ( );
FILL FILL_23_DFFSR_220 ( );
FILL FILL_24_DFFSR_220 ( );
FILL FILL_25_DFFSR_220 ( );
FILL FILL_26_DFFSR_220 ( );
FILL FILL_27_DFFSR_220 ( );
FILL FILL_28_DFFSR_220 ( );
FILL FILL_29_DFFSR_220 ( );
FILL FILL_30_DFFSR_220 ( );
FILL FILL_31_DFFSR_220 ( );
FILL FILL_32_DFFSR_220 ( );
FILL FILL_33_DFFSR_220 ( );
FILL FILL_34_DFFSR_220 ( );
FILL FILL_35_DFFSR_220 ( );
FILL FILL_36_DFFSR_220 ( );
FILL FILL_37_DFFSR_220 ( );
FILL FILL_38_DFFSR_220 ( );
FILL FILL_39_DFFSR_220 ( );
FILL FILL_40_DFFSR_220 ( );
FILL FILL_41_DFFSR_220 ( );
FILL FILL_42_DFFSR_220 ( );
FILL FILL_43_DFFSR_220 ( );
FILL FILL_44_DFFSR_220 ( );
FILL FILL_45_DFFSR_220 ( );
FILL FILL_46_DFFSR_220 ( );
FILL FILL_47_DFFSR_220 ( );
FILL FILL_48_DFFSR_220 ( );
FILL FILL_49_DFFSR_220 ( );
FILL FILL_50_DFFSR_220 ( );
FILL FILL_51_DFFSR_220 ( );
FILL FILL_0_DFFSR_227 ( );
FILL FILL_1_DFFSR_227 ( );
FILL FILL_2_DFFSR_227 ( );
FILL FILL_3_DFFSR_227 ( );
FILL FILL_4_DFFSR_227 ( );
FILL FILL_5_DFFSR_227 ( );
FILL FILL_6_DFFSR_227 ( );
FILL FILL_7_DFFSR_227 ( );
FILL FILL_8_DFFSR_227 ( );
FILL FILL_9_DFFSR_227 ( );
FILL FILL_10_DFFSR_227 ( );
FILL FILL_11_DFFSR_227 ( );
FILL FILL_12_DFFSR_227 ( );
FILL FILL_13_DFFSR_227 ( );
FILL FILL_14_DFFSR_227 ( );
FILL FILL_15_DFFSR_227 ( );
FILL FILL_16_DFFSR_227 ( );
FILL FILL_17_DFFSR_227 ( );
FILL FILL_18_DFFSR_227 ( );
FILL FILL_19_DFFSR_227 ( );
FILL FILL_20_DFFSR_227 ( );
FILL FILL_21_DFFSR_227 ( );
FILL FILL_22_DFFSR_227 ( );
FILL FILL_23_DFFSR_227 ( );
FILL FILL_24_DFFSR_227 ( );
FILL FILL_25_DFFSR_227 ( );
FILL FILL_26_DFFSR_227 ( );
FILL FILL_27_DFFSR_227 ( );
FILL FILL_28_DFFSR_227 ( );
FILL FILL_29_DFFSR_227 ( );
FILL FILL_30_DFFSR_227 ( );
FILL FILL_31_DFFSR_227 ( );
FILL FILL_32_DFFSR_227 ( );
FILL FILL_33_DFFSR_227 ( );
FILL FILL_34_DFFSR_227 ( );
FILL FILL_35_DFFSR_227 ( );
FILL FILL_36_DFFSR_227 ( );
FILL FILL_37_DFFSR_227 ( );
FILL FILL_38_DFFSR_227 ( );
FILL FILL_39_DFFSR_227 ( );
FILL FILL_40_DFFSR_227 ( );
FILL FILL_41_DFFSR_227 ( );
FILL FILL_42_DFFSR_227 ( );
FILL FILL_43_DFFSR_227 ( );
FILL FILL_44_DFFSR_227 ( );
FILL FILL_45_DFFSR_227 ( );
FILL FILL_46_DFFSR_227 ( );
FILL FILL_47_DFFSR_227 ( );
FILL FILL_48_DFFSR_227 ( );
FILL FILL_49_DFFSR_227 ( );
FILL FILL_50_DFFSR_227 ( );
FILL FILL_0_AOI22X1_11 ( );
FILL FILL_1_AOI22X1_11 ( );
FILL FILL_2_AOI22X1_11 ( );
FILL FILL_3_AOI22X1_11 ( );
FILL FILL_4_AOI22X1_11 ( );
FILL FILL_5_AOI22X1_11 ( );
FILL FILL_6_AOI22X1_11 ( );
FILL FILL_7_AOI22X1_11 ( );
FILL FILL_8_AOI22X1_11 ( );
FILL FILL_9_AOI22X1_11 ( );
FILL FILL_10_AOI22X1_11 ( );
FILL FILL_11_AOI22X1_11 ( );
FILL FILL_0_DFFSR_243 ( );
FILL FILL_1_DFFSR_243 ( );
FILL FILL_2_DFFSR_243 ( );
FILL FILL_3_DFFSR_243 ( );
FILL FILL_4_DFFSR_243 ( );
FILL FILL_5_DFFSR_243 ( );
FILL FILL_6_DFFSR_243 ( );
FILL FILL_7_DFFSR_243 ( );
FILL FILL_8_DFFSR_243 ( );
FILL FILL_9_DFFSR_243 ( );
FILL FILL_10_DFFSR_243 ( );
FILL FILL_11_DFFSR_243 ( );
FILL FILL_12_DFFSR_243 ( );
FILL FILL_13_DFFSR_243 ( );
FILL FILL_14_DFFSR_243 ( );
FILL FILL_15_DFFSR_243 ( );
FILL FILL_16_DFFSR_243 ( );
FILL FILL_17_DFFSR_243 ( );
FILL FILL_18_DFFSR_243 ( );
FILL FILL_19_DFFSR_243 ( );
FILL FILL_20_DFFSR_243 ( );
FILL FILL_21_DFFSR_243 ( );
FILL FILL_22_DFFSR_243 ( );
FILL FILL_23_DFFSR_243 ( );
FILL FILL_24_DFFSR_243 ( );
FILL FILL_25_DFFSR_243 ( );
FILL FILL_26_DFFSR_243 ( );
FILL FILL_27_DFFSR_243 ( );
FILL FILL_28_DFFSR_243 ( );
FILL FILL_29_DFFSR_243 ( );
FILL FILL_30_DFFSR_243 ( );
FILL FILL_31_DFFSR_243 ( );
FILL FILL_32_DFFSR_243 ( );
FILL FILL_33_DFFSR_243 ( );
FILL FILL_34_DFFSR_243 ( );
FILL FILL_35_DFFSR_243 ( );
FILL FILL_36_DFFSR_243 ( );
FILL FILL_37_DFFSR_243 ( );
FILL FILL_38_DFFSR_243 ( );
FILL FILL_39_DFFSR_243 ( );
FILL FILL_40_DFFSR_243 ( );
FILL FILL_41_DFFSR_243 ( );
FILL FILL_42_DFFSR_243 ( );
FILL FILL_43_DFFSR_243 ( );
FILL FILL_44_DFFSR_243 ( );
FILL FILL_45_DFFSR_243 ( );
FILL FILL_46_DFFSR_243 ( );
FILL FILL_47_DFFSR_243 ( );
FILL FILL_48_DFFSR_243 ( );
FILL FILL_49_DFFSR_243 ( );
FILL FILL_50_DFFSR_243 ( );
FILL FILL_0_NAND3X1_66 ( );
FILL FILL_1_NAND3X1_66 ( );
FILL FILL_2_NAND3X1_66 ( );
FILL FILL_3_NAND3X1_66 ( );
FILL FILL_4_NAND3X1_66 ( );
FILL FILL_5_NAND3X1_66 ( );
FILL FILL_6_NAND3X1_66 ( );
FILL FILL_7_NAND3X1_66 ( );
FILL FILL_8_NAND3X1_66 ( );
FILL FILL_0_NAND2X1_41 ( );
FILL FILL_1_NAND2X1_41 ( );
FILL FILL_2_NAND2X1_41 ( );
FILL FILL_3_NAND2X1_41 ( );
FILL FILL_4_NAND2X1_41 ( );
FILL FILL_5_NAND2X1_41 ( );
FILL FILL_6_NAND2X1_41 ( );
FILL FILL_0_DFFSR_251 ( );
FILL FILL_1_DFFSR_251 ( );
FILL FILL_2_DFFSR_251 ( );
FILL FILL_3_DFFSR_251 ( );
FILL FILL_4_DFFSR_251 ( );
FILL FILL_5_DFFSR_251 ( );
FILL FILL_6_DFFSR_251 ( );
FILL FILL_7_DFFSR_251 ( );
FILL FILL_8_DFFSR_251 ( );
FILL FILL_9_DFFSR_251 ( );
FILL FILL_10_DFFSR_251 ( );
FILL FILL_11_DFFSR_251 ( );
FILL FILL_12_DFFSR_251 ( );
FILL FILL_13_DFFSR_251 ( );
FILL FILL_14_DFFSR_251 ( );
FILL FILL_15_DFFSR_251 ( );
FILL FILL_16_DFFSR_251 ( );
FILL FILL_17_DFFSR_251 ( );
FILL FILL_18_DFFSR_251 ( );
FILL FILL_19_DFFSR_251 ( );
FILL FILL_20_DFFSR_251 ( );
FILL FILL_21_DFFSR_251 ( );
FILL FILL_22_DFFSR_251 ( );
FILL FILL_23_DFFSR_251 ( );
FILL FILL_24_DFFSR_251 ( );
FILL FILL_25_DFFSR_251 ( );
FILL FILL_26_DFFSR_251 ( );
FILL FILL_27_DFFSR_251 ( );
FILL FILL_28_DFFSR_251 ( );
FILL FILL_29_DFFSR_251 ( );
FILL FILL_30_DFFSR_251 ( );
FILL FILL_31_DFFSR_251 ( );
FILL FILL_32_DFFSR_251 ( );
FILL FILL_33_DFFSR_251 ( );
FILL FILL_34_DFFSR_251 ( );
FILL FILL_35_DFFSR_251 ( );
FILL FILL_36_DFFSR_251 ( );
FILL FILL_37_DFFSR_251 ( );
FILL FILL_38_DFFSR_251 ( );
FILL FILL_39_DFFSR_251 ( );
FILL FILL_40_DFFSR_251 ( );
FILL FILL_41_DFFSR_251 ( );
FILL FILL_42_DFFSR_251 ( );
FILL FILL_43_DFFSR_251 ( );
FILL FILL_44_DFFSR_251 ( );
FILL FILL_45_DFFSR_251 ( );
FILL FILL_46_DFFSR_251 ( );
FILL FILL_47_DFFSR_251 ( );
FILL FILL_48_DFFSR_251 ( );
FILL FILL_49_DFFSR_251 ( );
FILL FILL_50_DFFSR_251 ( );
FILL FILL_51_DFFSR_251 ( );
FILL FILL_0_INVX1_65 ( );
FILL FILL_1_INVX1_65 ( );
FILL FILL_2_INVX1_65 ( );
FILL FILL_3_INVX1_65 ( );
FILL FILL_4_INVX1_65 ( );
FILL FILL_0_NAND3X1_70 ( );
FILL FILL_1_NAND3X1_70 ( );
FILL FILL_2_NAND3X1_70 ( );
FILL FILL_3_NAND3X1_70 ( );
FILL FILL_4_NAND3X1_70 ( );
FILL FILL_5_NAND3X1_70 ( );
FILL FILL_6_NAND3X1_70 ( );
FILL FILL_7_NAND3X1_70 ( );
FILL FILL_8_NAND3X1_70 ( );
FILL FILL_9_NAND3X1_70 ( );
FILL FILL_0_INVX1_104 ( );
FILL FILL_1_INVX1_104 ( );
FILL FILL_2_INVX1_104 ( );
FILL FILL_3_INVX1_104 ( );
FILL FILL_0_INVX1_105 ( );
FILL FILL_1_INVX1_105 ( );
FILL FILL_2_INVX1_105 ( );
FILL FILL_3_INVX1_105 ( );
FILL FILL_4_INVX1_105 ( );
FILL FILL_0_INVX1_117 ( );
FILL FILL_1_INVX1_117 ( );
FILL FILL_2_INVX1_117 ( );
FILL FILL_3_INVX1_117 ( );
FILL FILL_4_INVX1_117 ( );
FILL FILL_0_DFFSR_224 ( );
FILL FILL_1_DFFSR_224 ( );
FILL FILL_2_DFFSR_224 ( );
FILL FILL_3_DFFSR_224 ( );
FILL FILL_4_DFFSR_224 ( );
FILL FILL_5_DFFSR_224 ( );
FILL FILL_6_DFFSR_224 ( );
FILL FILL_7_DFFSR_224 ( );
FILL FILL_8_DFFSR_224 ( );
FILL FILL_9_DFFSR_224 ( );
FILL FILL_10_DFFSR_224 ( );
FILL FILL_11_DFFSR_224 ( );
FILL FILL_12_DFFSR_224 ( );
FILL FILL_13_DFFSR_224 ( );
FILL FILL_14_DFFSR_224 ( );
FILL FILL_15_DFFSR_224 ( );
FILL FILL_16_DFFSR_224 ( );
FILL FILL_17_DFFSR_224 ( );
FILL FILL_18_DFFSR_224 ( );
FILL FILL_19_DFFSR_224 ( );
FILL FILL_20_DFFSR_224 ( );
FILL FILL_21_DFFSR_224 ( );
FILL FILL_22_DFFSR_224 ( );
FILL FILL_23_DFFSR_224 ( );
FILL FILL_24_DFFSR_224 ( );
FILL FILL_25_DFFSR_224 ( );
FILL FILL_26_DFFSR_224 ( );
FILL FILL_27_DFFSR_224 ( );
FILL FILL_28_DFFSR_224 ( );
FILL FILL_29_DFFSR_224 ( );
FILL FILL_30_DFFSR_224 ( );
FILL FILL_31_DFFSR_224 ( );
FILL FILL_32_DFFSR_224 ( );
FILL FILL_33_DFFSR_224 ( );
FILL FILL_34_DFFSR_224 ( );
FILL FILL_35_DFFSR_224 ( );
FILL FILL_36_DFFSR_224 ( );
FILL FILL_37_DFFSR_224 ( );
FILL FILL_38_DFFSR_224 ( );
FILL FILL_39_DFFSR_224 ( );
FILL FILL_40_DFFSR_224 ( );
FILL FILL_41_DFFSR_224 ( );
FILL FILL_42_DFFSR_224 ( );
FILL FILL_43_DFFSR_224 ( );
FILL FILL_44_DFFSR_224 ( );
FILL FILL_45_DFFSR_224 ( );
FILL FILL_46_DFFSR_224 ( );
FILL FILL_47_DFFSR_224 ( );
FILL FILL_48_DFFSR_224 ( );
FILL FILL_49_DFFSR_224 ( );
FILL FILL_50_DFFSR_224 ( );
FILL FILL_0_OAI21X1_53 ( );
FILL FILL_1_OAI21X1_53 ( );
FILL FILL_2_OAI21X1_53 ( );
FILL FILL_3_OAI21X1_53 ( );
FILL FILL_4_OAI21X1_53 ( );
FILL FILL_5_OAI21X1_53 ( );
FILL FILL_6_OAI21X1_53 ( );
FILL FILL_7_OAI21X1_53 ( );
FILL FILL_8_OAI21X1_53 ( );
FILL FILL_0_DFFSR_278 ( );
FILL FILL_1_DFFSR_278 ( );
FILL FILL_2_DFFSR_278 ( );
FILL FILL_3_DFFSR_278 ( );
FILL FILL_4_DFFSR_278 ( );
FILL FILL_5_DFFSR_278 ( );
FILL FILL_6_DFFSR_278 ( );
FILL FILL_7_DFFSR_278 ( );
FILL FILL_8_DFFSR_278 ( );
FILL FILL_9_DFFSR_278 ( );
FILL FILL_10_DFFSR_278 ( );
FILL FILL_11_DFFSR_278 ( );
FILL FILL_12_DFFSR_278 ( );
FILL FILL_13_DFFSR_278 ( );
FILL FILL_14_DFFSR_278 ( );
FILL FILL_15_DFFSR_278 ( );
FILL FILL_16_DFFSR_278 ( );
FILL FILL_17_DFFSR_278 ( );
FILL FILL_18_DFFSR_278 ( );
FILL FILL_19_DFFSR_278 ( );
FILL FILL_20_DFFSR_278 ( );
FILL FILL_21_DFFSR_278 ( );
FILL FILL_22_DFFSR_278 ( );
FILL FILL_23_DFFSR_278 ( );
FILL FILL_24_DFFSR_278 ( );
FILL FILL_25_DFFSR_278 ( );
FILL FILL_26_DFFSR_278 ( );
FILL FILL_27_DFFSR_278 ( );
FILL FILL_28_DFFSR_278 ( );
FILL FILL_29_DFFSR_278 ( );
FILL FILL_30_DFFSR_278 ( );
FILL FILL_31_DFFSR_278 ( );
FILL FILL_32_DFFSR_278 ( );
FILL FILL_33_DFFSR_278 ( );
FILL FILL_34_DFFSR_278 ( );
FILL FILL_35_DFFSR_278 ( );
FILL FILL_36_DFFSR_278 ( );
FILL FILL_37_DFFSR_278 ( );
FILL FILL_38_DFFSR_278 ( );
FILL FILL_39_DFFSR_278 ( );
FILL FILL_40_DFFSR_278 ( );
FILL FILL_41_DFFSR_278 ( );
FILL FILL_42_DFFSR_278 ( );
FILL FILL_43_DFFSR_278 ( );
FILL FILL_44_DFFSR_278 ( );
FILL FILL_45_DFFSR_278 ( );
FILL FILL_46_DFFSR_278 ( );
FILL FILL_47_DFFSR_278 ( );
FILL FILL_48_DFFSR_278 ( );
FILL FILL_49_DFFSR_278 ( );
FILL FILL_50_DFFSR_278 ( );
FILL FILL_51_DFFSR_278 ( );
FILL FILL_0_AOI21X1_9 ( );
FILL FILL_1_AOI21X1_9 ( );
FILL FILL_2_AOI21X1_9 ( );
FILL FILL_3_AOI21X1_9 ( );
FILL FILL_4_AOI21X1_9 ( );
FILL FILL_5_AOI21X1_9 ( );
FILL FILL_6_AOI21X1_9 ( );
FILL FILL_7_AOI21X1_9 ( );
FILL FILL_8_AOI21X1_9 ( );
FILL FILL_0_NAND3X1_153 ( );
FILL FILL_1_NAND3X1_153 ( );
FILL FILL_2_NAND3X1_153 ( );
FILL FILL_3_NAND3X1_153 ( );
FILL FILL_4_NAND3X1_153 ( );
FILL FILL_5_NAND3X1_153 ( );
FILL FILL_6_NAND3X1_153 ( );
FILL FILL_7_NAND3X1_153 ( );
FILL FILL_8_NAND3X1_153 ( );
FILL FILL_0_NAND2X1_79 ( );
FILL FILL_1_NAND2X1_79 ( );
FILL FILL_2_NAND2X1_79 ( );
FILL FILL_3_NAND2X1_79 ( );
FILL FILL_4_NAND2X1_79 ( );
FILL FILL_5_NAND2X1_79 ( );
FILL FILL_6_NAND2X1_79 ( );
FILL FILL_0_NAND2X1_65 ( );
FILL FILL_1_NAND2X1_65 ( );
FILL FILL_2_NAND2X1_65 ( );
FILL FILL_3_NAND2X1_65 ( );
FILL FILL_4_NAND2X1_65 ( );
FILL FILL_5_NAND2X1_65 ( );
FILL FILL_6_NAND2X1_65 ( );
FILL FILL_0_NAND2X1_132 ( );
FILL FILL_1_NAND2X1_132 ( );
FILL FILL_2_NAND2X1_132 ( );
FILL FILL_3_NAND2X1_132 ( );
FILL FILL_4_NAND2X1_132 ( );
FILL FILL_5_NAND2X1_132 ( );
FILL FILL_6_NAND2X1_132 ( );
FILL FILL_0_OAI21X1_28 ( );
FILL FILL_1_OAI21X1_28 ( );
FILL FILL_2_OAI21X1_28 ( );
FILL FILL_3_OAI21X1_28 ( );
FILL FILL_4_OAI21X1_28 ( );
FILL FILL_5_OAI21X1_28 ( );
FILL FILL_6_OAI21X1_28 ( );
FILL FILL_7_OAI21X1_28 ( );
FILL FILL_8_OAI21X1_28 ( );
FILL FILL_9_OAI21X1_28 ( );
FILL FILL_0_BUFX2_52 ( );
FILL FILL_1_BUFX2_52 ( );
FILL FILL_2_BUFX2_52 ( );
FILL FILL_3_BUFX2_52 ( );
FILL FILL_4_BUFX2_52 ( );
FILL FILL_5_BUFX2_52 ( );
FILL FILL_6_BUFX2_52 ( );
FILL FILL_0_INVX1_192 ( );
FILL FILL_1_INVX1_192 ( );
FILL FILL_2_INVX1_192 ( );
FILL FILL_3_INVX1_192 ( );
FILL FILL_0_NAND2X1_145 ( );
FILL FILL_1_NAND2X1_145 ( );
FILL FILL_2_NAND2X1_145 ( );
FILL FILL_3_NAND2X1_145 ( );
FILL FILL_4_NAND2X1_145 ( );
FILL FILL_5_NAND2X1_145 ( );
FILL FILL_6_NAND2X1_145 ( );
FILL FILL_0_DFFSR_142 ( );
FILL FILL_1_DFFSR_142 ( );
FILL FILL_2_DFFSR_142 ( );
FILL FILL_3_DFFSR_142 ( );
FILL FILL_4_DFFSR_142 ( );
FILL FILL_5_DFFSR_142 ( );
FILL FILL_6_DFFSR_142 ( );
FILL FILL_7_DFFSR_142 ( );
FILL FILL_8_DFFSR_142 ( );
FILL FILL_9_DFFSR_142 ( );
FILL FILL_10_DFFSR_142 ( );
FILL FILL_11_DFFSR_142 ( );
FILL FILL_12_DFFSR_142 ( );
FILL FILL_13_DFFSR_142 ( );
FILL FILL_14_DFFSR_142 ( );
FILL FILL_15_DFFSR_142 ( );
FILL FILL_16_DFFSR_142 ( );
FILL FILL_17_DFFSR_142 ( );
FILL FILL_18_DFFSR_142 ( );
FILL FILL_19_DFFSR_142 ( );
FILL FILL_20_DFFSR_142 ( );
FILL FILL_21_DFFSR_142 ( );
FILL FILL_22_DFFSR_142 ( );
FILL FILL_23_DFFSR_142 ( );
FILL FILL_24_DFFSR_142 ( );
FILL FILL_25_DFFSR_142 ( );
FILL FILL_26_DFFSR_142 ( );
FILL FILL_27_DFFSR_142 ( );
FILL FILL_28_DFFSR_142 ( );
FILL FILL_29_DFFSR_142 ( );
FILL FILL_30_DFFSR_142 ( );
FILL FILL_31_DFFSR_142 ( );
FILL FILL_32_DFFSR_142 ( );
FILL FILL_33_DFFSR_142 ( );
FILL FILL_34_DFFSR_142 ( );
FILL FILL_35_DFFSR_142 ( );
FILL FILL_36_DFFSR_142 ( );
FILL FILL_37_DFFSR_142 ( );
FILL FILL_38_DFFSR_142 ( );
FILL FILL_39_DFFSR_142 ( );
FILL FILL_40_DFFSR_142 ( );
FILL FILL_41_DFFSR_142 ( );
FILL FILL_42_DFFSR_142 ( );
FILL FILL_43_DFFSR_142 ( );
FILL FILL_44_DFFSR_142 ( );
FILL FILL_45_DFFSR_142 ( );
FILL FILL_46_DFFSR_142 ( );
FILL FILL_47_DFFSR_142 ( );
FILL FILL_48_DFFSR_142 ( );
FILL FILL_49_DFFSR_142 ( );
FILL FILL_50_DFFSR_142 ( );
FILL FILL_0_CLKBUF1_21 ( );
FILL FILL_1_CLKBUF1_21 ( );
FILL FILL_2_CLKBUF1_21 ( );
FILL FILL_3_CLKBUF1_21 ( );
FILL FILL_4_CLKBUF1_21 ( );
FILL FILL_5_CLKBUF1_21 ( );
FILL FILL_6_CLKBUF1_21 ( );
FILL FILL_7_CLKBUF1_21 ( );
FILL FILL_8_CLKBUF1_21 ( );
FILL FILL_9_CLKBUF1_21 ( );
FILL FILL_10_CLKBUF1_21 ( );
FILL FILL_11_CLKBUF1_21 ( );
FILL FILL_12_CLKBUF1_21 ( );
FILL FILL_13_CLKBUF1_21 ( );
FILL FILL_14_CLKBUF1_21 ( );
FILL FILL_15_CLKBUF1_21 ( );
FILL FILL_16_CLKBUF1_21 ( );
FILL FILL_17_CLKBUF1_21 ( );
FILL FILL_18_CLKBUF1_21 ( );
FILL FILL_19_CLKBUF1_21 ( );
FILL FILL_20_CLKBUF1_21 ( );
FILL FILL_0_DFFSR_196 ( );
FILL FILL_1_DFFSR_196 ( );
FILL FILL_2_DFFSR_196 ( );
FILL FILL_3_DFFSR_196 ( );
FILL FILL_4_DFFSR_196 ( );
FILL FILL_5_DFFSR_196 ( );
FILL FILL_6_DFFSR_196 ( );
FILL FILL_7_DFFSR_196 ( );
FILL FILL_8_DFFSR_196 ( );
FILL FILL_9_DFFSR_196 ( );
FILL FILL_10_DFFSR_196 ( );
FILL FILL_11_DFFSR_196 ( );
FILL FILL_12_DFFSR_196 ( );
FILL FILL_13_DFFSR_196 ( );
FILL FILL_14_DFFSR_196 ( );
FILL FILL_15_DFFSR_196 ( );
FILL FILL_16_DFFSR_196 ( );
FILL FILL_17_DFFSR_196 ( );
FILL FILL_18_DFFSR_196 ( );
FILL FILL_19_DFFSR_196 ( );
FILL FILL_20_DFFSR_196 ( );
FILL FILL_21_DFFSR_196 ( );
FILL FILL_22_DFFSR_196 ( );
FILL FILL_23_DFFSR_196 ( );
FILL FILL_24_DFFSR_196 ( );
FILL FILL_25_DFFSR_196 ( );
FILL FILL_26_DFFSR_196 ( );
FILL FILL_27_DFFSR_196 ( );
FILL FILL_28_DFFSR_196 ( );
FILL FILL_29_DFFSR_196 ( );
FILL FILL_30_DFFSR_196 ( );
FILL FILL_31_DFFSR_196 ( );
FILL FILL_32_DFFSR_196 ( );
FILL FILL_33_DFFSR_196 ( );
FILL FILL_34_DFFSR_196 ( );
FILL FILL_35_DFFSR_196 ( );
FILL FILL_36_DFFSR_196 ( );
FILL FILL_37_DFFSR_196 ( );
FILL FILL_38_DFFSR_196 ( );
FILL FILL_39_DFFSR_196 ( );
FILL FILL_40_DFFSR_196 ( );
FILL FILL_41_DFFSR_196 ( );
FILL FILL_42_DFFSR_196 ( );
FILL FILL_43_DFFSR_196 ( );
FILL FILL_44_DFFSR_196 ( );
FILL FILL_45_DFFSR_196 ( );
FILL FILL_46_DFFSR_196 ( );
FILL FILL_47_DFFSR_196 ( );
FILL FILL_48_DFFSR_196 ( );
FILL FILL_49_DFFSR_196 ( );
FILL FILL_50_DFFSR_196 ( );
FILL FILL_51_DFFSR_196 ( );
FILL FILL_0_NAND3X1_110 ( );
FILL FILL_1_NAND3X1_110 ( );
FILL FILL_2_NAND3X1_110 ( );
FILL FILL_3_NAND3X1_110 ( );
FILL FILL_4_NAND3X1_110 ( );
FILL FILL_5_NAND3X1_110 ( );
FILL FILL_6_NAND3X1_110 ( );
FILL FILL_7_NAND3X1_110 ( );
FILL FILL_8_NAND3X1_110 ( );
FILL FILL_0_NAND3X1_111 ( );
FILL FILL_1_NAND3X1_111 ( );
FILL FILL_2_NAND3X1_111 ( );
FILL FILL_3_NAND3X1_111 ( );
FILL FILL_4_NAND3X1_111 ( );
FILL FILL_5_NAND3X1_111 ( );
FILL FILL_6_NAND3X1_111 ( );
FILL FILL_7_NAND3X1_111 ( );
FILL FILL_8_NAND3X1_111 ( );
FILL FILL_0_NAND3X1_109 ( );
FILL FILL_1_NAND3X1_109 ( );
FILL FILL_2_NAND3X1_109 ( );
FILL FILL_3_NAND3X1_109 ( );
FILL FILL_4_NAND3X1_109 ( );
FILL FILL_5_NAND3X1_109 ( );
FILL FILL_6_NAND3X1_109 ( );
FILL FILL_7_NAND3X1_109 ( );
FILL FILL_8_NAND3X1_109 ( );
FILL FILL_0_DFFSR_129 ( );
FILL FILL_1_DFFSR_129 ( );
FILL FILL_2_DFFSR_129 ( );
FILL FILL_3_DFFSR_129 ( );
FILL FILL_4_DFFSR_129 ( );
FILL FILL_5_DFFSR_129 ( );
FILL FILL_6_DFFSR_129 ( );
FILL FILL_7_DFFSR_129 ( );
FILL FILL_8_DFFSR_129 ( );
FILL FILL_9_DFFSR_129 ( );
FILL FILL_10_DFFSR_129 ( );
FILL FILL_11_DFFSR_129 ( );
FILL FILL_12_DFFSR_129 ( );
FILL FILL_13_DFFSR_129 ( );
FILL FILL_14_DFFSR_129 ( );
FILL FILL_15_DFFSR_129 ( );
FILL FILL_16_DFFSR_129 ( );
FILL FILL_17_DFFSR_129 ( );
FILL FILL_18_DFFSR_129 ( );
FILL FILL_19_DFFSR_129 ( );
FILL FILL_20_DFFSR_129 ( );
FILL FILL_21_DFFSR_129 ( );
FILL FILL_22_DFFSR_129 ( );
FILL FILL_23_DFFSR_129 ( );
FILL FILL_24_DFFSR_129 ( );
FILL FILL_25_DFFSR_129 ( );
FILL FILL_26_DFFSR_129 ( );
FILL FILL_27_DFFSR_129 ( );
FILL FILL_28_DFFSR_129 ( );
FILL FILL_29_DFFSR_129 ( );
FILL FILL_30_DFFSR_129 ( );
FILL FILL_31_DFFSR_129 ( );
FILL FILL_32_DFFSR_129 ( );
FILL FILL_33_DFFSR_129 ( );
FILL FILL_34_DFFSR_129 ( );
FILL FILL_35_DFFSR_129 ( );
FILL FILL_36_DFFSR_129 ( );
FILL FILL_37_DFFSR_129 ( );
FILL FILL_38_DFFSR_129 ( );
FILL FILL_39_DFFSR_129 ( );
FILL FILL_40_DFFSR_129 ( );
FILL FILL_41_DFFSR_129 ( );
FILL FILL_42_DFFSR_129 ( );
FILL FILL_43_DFFSR_129 ( );
FILL FILL_44_DFFSR_129 ( );
FILL FILL_45_DFFSR_129 ( );
FILL FILL_46_DFFSR_129 ( );
FILL FILL_47_DFFSR_129 ( );
FILL FILL_48_DFFSR_129 ( );
FILL FILL_49_DFFSR_129 ( );
FILL FILL_50_DFFSR_129 ( );
FILL FILL_0_NAND3X1_67 ( );
FILL FILL_1_NAND3X1_67 ( );
FILL FILL_2_NAND3X1_67 ( );
FILL FILL_3_NAND3X1_67 ( );
FILL FILL_4_NAND3X1_67 ( );
FILL FILL_5_NAND3X1_67 ( );
FILL FILL_6_NAND3X1_67 ( );
FILL FILL_7_NAND3X1_67 ( );
FILL FILL_8_NAND3X1_67 ( );
FILL FILL_0_BUFX2_23 ( );
FILL FILL_1_BUFX2_23 ( );
FILL FILL_2_BUFX2_23 ( );
FILL FILL_3_BUFX2_23 ( );
FILL FILL_4_BUFX2_23 ( );
FILL FILL_5_BUFX2_23 ( );
FILL FILL_6_BUFX2_23 ( );
FILL FILL_0_BUFX2_92 ( );
FILL FILL_1_BUFX2_92 ( );
FILL FILL_2_BUFX2_92 ( );
FILL FILL_3_BUFX2_92 ( );
FILL FILL_4_BUFX2_92 ( );
FILL FILL_5_BUFX2_92 ( );
FILL FILL_6_BUFX2_92 ( );
FILL FILL_0_INVX1_82 ( );
FILL FILL_1_INVX1_82 ( );
FILL FILL_2_INVX1_82 ( );
FILL FILL_3_INVX1_82 ( );
FILL FILL_4_INVX1_82 ( );
FILL FILL_0_NAND3X1_83 ( );
FILL FILL_1_NAND3X1_83 ( );
FILL FILL_2_NAND3X1_83 ( );
FILL FILL_3_NAND3X1_83 ( );
FILL FILL_4_NAND3X1_83 ( );
FILL FILL_5_NAND3X1_83 ( );
FILL FILL_6_NAND3X1_83 ( );
FILL FILL_7_NAND3X1_83 ( );
FILL FILL_8_NAND3X1_83 ( );
FILL FILL_0_BUFX2_24 ( );
FILL FILL_1_BUFX2_24 ( );
FILL FILL_2_BUFX2_24 ( );
FILL FILL_3_BUFX2_24 ( );
FILL FILL_4_BUFX2_24 ( );
FILL FILL_5_BUFX2_24 ( );
FILL FILL_6_BUFX2_24 ( );
FILL FILL_0_DFFSR_157 ( );
FILL FILL_1_DFFSR_157 ( );
FILL FILL_2_DFFSR_157 ( );
FILL FILL_3_DFFSR_157 ( );
FILL FILL_4_DFFSR_157 ( );
FILL FILL_5_DFFSR_157 ( );
FILL FILL_6_DFFSR_157 ( );
FILL FILL_7_DFFSR_157 ( );
FILL FILL_8_DFFSR_157 ( );
FILL FILL_9_DFFSR_157 ( );
FILL FILL_10_DFFSR_157 ( );
FILL FILL_11_DFFSR_157 ( );
FILL FILL_12_DFFSR_157 ( );
FILL FILL_13_DFFSR_157 ( );
FILL FILL_14_DFFSR_157 ( );
FILL FILL_15_DFFSR_157 ( );
FILL FILL_16_DFFSR_157 ( );
FILL FILL_17_DFFSR_157 ( );
FILL FILL_18_DFFSR_157 ( );
FILL FILL_19_DFFSR_157 ( );
FILL FILL_20_DFFSR_157 ( );
FILL FILL_21_DFFSR_157 ( );
FILL FILL_22_DFFSR_157 ( );
FILL FILL_23_DFFSR_157 ( );
FILL FILL_24_DFFSR_157 ( );
FILL FILL_25_DFFSR_157 ( );
FILL FILL_26_DFFSR_157 ( );
FILL FILL_27_DFFSR_157 ( );
FILL FILL_28_DFFSR_157 ( );
FILL FILL_29_DFFSR_157 ( );
FILL FILL_30_DFFSR_157 ( );
FILL FILL_31_DFFSR_157 ( );
FILL FILL_32_DFFSR_157 ( );
FILL FILL_33_DFFSR_157 ( );
FILL FILL_34_DFFSR_157 ( );
FILL FILL_35_DFFSR_157 ( );
FILL FILL_36_DFFSR_157 ( );
FILL FILL_37_DFFSR_157 ( );
FILL FILL_38_DFFSR_157 ( );
FILL FILL_39_DFFSR_157 ( );
FILL FILL_40_DFFSR_157 ( );
FILL FILL_41_DFFSR_157 ( );
FILL FILL_42_DFFSR_157 ( );
FILL FILL_43_DFFSR_157 ( );
FILL FILL_44_DFFSR_157 ( );
FILL FILL_45_DFFSR_157 ( );
FILL FILL_46_DFFSR_157 ( );
FILL FILL_47_DFFSR_157 ( );
FILL FILL_48_DFFSR_157 ( );
FILL FILL_49_DFFSR_157 ( );
FILL FILL_50_DFFSR_157 ( );
FILL FILL_0_DFFSR_151 ( );
FILL FILL_1_DFFSR_151 ( );
FILL FILL_2_DFFSR_151 ( );
FILL FILL_3_DFFSR_151 ( );
FILL FILL_4_DFFSR_151 ( );
FILL FILL_5_DFFSR_151 ( );
FILL FILL_6_DFFSR_151 ( );
FILL FILL_7_DFFSR_151 ( );
FILL FILL_8_DFFSR_151 ( );
FILL FILL_9_DFFSR_151 ( );
FILL FILL_10_DFFSR_151 ( );
FILL FILL_11_DFFSR_151 ( );
FILL FILL_12_DFFSR_151 ( );
FILL FILL_13_DFFSR_151 ( );
FILL FILL_14_DFFSR_151 ( );
FILL FILL_15_DFFSR_151 ( );
FILL FILL_16_DFFSR_151 ( );
FILL FILL_17_DFFSR_151 ( );
FILL FILL_18_DFFSR_151 ( );
FILL FILL_19_DFFSR_151 ( );
FILL FILL_20_DFFSR_151 ( );
FILL FILL_21_DFFSR_151 ( );
FILL FILL_22_DFFSR_151 ( );
FILL FILL_23_DFFSR_151 ( );
FILL FILL_24_DFFSR_151 ( );
FILL FILL_25_DFFSR_151 ( );
FILL FILL_26_DFFSR_151 ( );
FILL FILL_27_DFFSR_151 ( );
FILL FILL_28_DFFSR_151 ( );
FILL FILL_29_DFFSR_151 ( );
FILL FILL_30_DFFSR_151 ( );
FILL FILL_31_DFFSR_151 ( );
FILL FILL_32_DFFSR_151 ( );
FILL FILL_33_DFFSR_151 ( );
FILL FILL_34_DFFSR_151 ( );
FILL FILL_35_DFFSR_151 ( );
FILL FILL_36_DFFSR_151 ( );
FILL FILL_37_DFFSR_151 ( );
FILL FILL_38_DFFSR_151 ( );
FILL FILL_39_DFFSR_151 ( );
FILL FILL_40_DFFSR_151 ( );
FILL FILL_41_DFFSR_151 ( );
FILL FILL_42_DFFSR_151 ( );
FILL FILL_43_DFFSR_151 ( );
FILL FILL_44_DFFSR_151 ( );
FILL FILL_45_DFFSR_151 ( );
FILL FILL_46_DFFSR_151 ( );
FILL FILL_47_DFFSR_151 ( );
FILL FILL_48_DFFSR_151 ( );
FILL FILL_49_DFFSR_151 ( );
FILL FILL_50_DFFSR_151 ( );
FILL FILL_0_OAI21X1_54 ( );
FILL FILL_1_OAI21X1_54 ( );
FILL FILL_2_OAI21X1_54 ( );
FILL FILL_3_OAI21X1_54 ( );
FILL FILL_4_OAI21X1_54 ( );
FILL FILL_5_OAI21X1_54 ( );
FILL FILL_6_OAI21X1_54 ( );
FILL FILL_7_OAI21X1_54 ( );
FILL FILL_8_OAI21X1_54 ( );
FILL FILL_9_OAI21X1_54 ( );
FILL FILL_0_OAI21X1_52 ( );
FILL FILL_1_OAI21X1_52 ( );
FILL FILL_2_OAI21X1_52 ( );
FILL FILL_3_OAI21X1_52 ( );
FILL FILL_4_OAI21X1_52 ( );
FILL FILL_5_OAI21X1_52 ( );
FILL FILL_6_OAI21X1_52 ( );
FILL FILL_7_OAI21X1_52 ( );
FILL FILL_8_OAI21X1_52 ( );
FILL FILL_9_OAI21X1_52 ( );
FILL FILL_0_AOI21X1_33 ( );
FILL FILL_1_AOI21X1_33 ( );
FILL FILL_2_AOI21X1_33 ( );
FILL FILL_3_AOI21X1_33 ( );
FILL FILL_4_AOI21X1_33 ( );
FILL FILL_5_AOI21X1_33 ( );
FILL FILL_6_AOI21X1_33 ( );
FILL FILL_7_AOI21X1_33 ( );
FILL FILL_8_AOI21X1_33 ( );
FILL FILL_0_OAI21X1_106 ( );
FILL FILL_1_OAI21X1_106 ( );
FILL FILL_2_OAI21X1_106 ( );
FILL FILL_3_OAI21X1_106 ( );
FILL FILL_4_OAI21X1_106 ( );
FILL FILL_5_OAI21X1_106 ( );
FILL FILL_6_OAI21X1_106 ( );
FILL FILL_7_OAI21X1_106 ( );
FILL FILL_8_OAI21X1_106 ( );
FILL FILL_0_NAND3X1_193 ( );
FILL FILL_1_NAND3X1_193 ( );
FILL FILL_2_NAND3X1_193 ( );
FILL FILL_3_NAND3X1_193 ( );
FILL FILL_4_NAND3X1_193 ( );
FILL FILL_5_NAND3X1_193 ( );
FILL FILL_6_NAND3X1_193 ( );
FILL FILL_7_NAND3X1_193 ( );
FILL FILL_8_NAND3X1_193 ( );
FILL FILL_0_NAND3X1_167 ( );
FILL FILL_1_NAND3X1_167 ( );
FILL FILL_2_NAND3X1_167 ( );
FILL FILL_3_NAND3X1_167 ( );
FILL FILL_4_NAND3X1_167 ( );
FILL FILL_5_NAND3X1_167 ( );
FILL FILL_6_NAND3X1_167 ( );
FILL FILL_7_NAND3X1_167 ( );
FILL FILL_8_NAND3X1_167 ( );
FILL FILL_0_XOR2X1_1 ( );
FILL FILL_1_XOR2X1_1 ( );
FILL FILL_2_XOR2X1_1 ( );
FILL FILL_3_XOR2X1_1 ( );
FILL FILL_4_XOR2X1_1 ( );
FILL FILL_5_XOR2X1_1 ( );
FILL FILL_6_XOR2X1_1 ( );
FILL FILL_7_XOR2X1_1 ( );
FILL FILL_8_XOR2X1_1 ( );
FILL FILL_9_XOR2X1_1 ( );
FILL FILL_10_XOR2X1_1 ( );
FILL FILL_11_XOR2X1_1 ( );
FILL FILL_12_XOR2X1_1 ( );
FILL FILL_13_XOR2X1_1 ( );
FILL FILL_14_XOR2X1_1 ( );
FILL FILL_15_XOR2X1_1 ( );
FILL FILL_16_XOR2X1_1 ( );
FILL FILL_0_NAND3X1_168 ( );
FILL FILL_1_NAND3X1_168 ( );
FILL FILL_2_NAND3X1_168 ( );
FILL FILL_3_NAND3X1_168 ( );
FILL FILL_4_NAND3X1_168 ( );
FILL FILL_5_NAND3X1_168 ( );
FILL FILL_6_NAND3X1_168 ( );
FILL FILL_7_NAND3X1_168 ( );
FILL FILL_8_NAND3X1_168 ( );
FILL FILL_0_INVX1_154 ( );
FILL FILL_1_INVX1_154 ( );
FILL FILL_2_INVX1_154 ( );
FILL FILL_3_INVX1_154 ( );
FILL FILL_4_INVX1_154 ( );
FILL FILL_0_NAND2X1_80 ( );
FILL FILL_1_NAND2X1_80 ( );
FILL FILL_2_NAND2X1_80 ( );
FILL FILL_3_NAND2X1_80 ( );
FILL FILL_4_NAND2X1_80 ( );
FILL FILL_5_NAND2X1_80 ( );
FILL FILL_6_NAND2X1_80 ( );
FILL FILL_0_NAND3X1_169 ( );
FILL FILL_1_NAND3X1_169 ( );
FILL FILL_2_NAND3X1_169 ( );
FILL FILL_3_NAND3X1_169 ( );
FILL FILL_4_NAND3X1_169 ( );
FILL FILL_5_NAND3X1_169 ( );
FILL FILL_6_NAND3X1_169 ( );
FILL FILL_7_NAND3X1_169 ( );
FILL FILL_8_NAND3X1_169 ( );
FILL FILL_0_NAND3X1_170 ( );
FILL FILL_1_NAND3X1_170 ( );
FILL FILL_2_NAND3X1_170 ( );
FILL FILL_3_NAND3X1_170 ( );
FILL FILL_4_NAND3X1_170 ( );
FILL FILL_5_NAND3X1_170 ( );
FILL FILL_6_NAND3X1_170 ( );
FILL FILL_7_NAND3X1_170 ( );
FILL FILL_8_NAND3X1_170 ( );
FILL FILL_0_DFFSR_267 ( );
FILL FILL_1_DFFSR_267 ( );
FILL FILL_2_DFFSR_267 ( );
FILL FILL_3_DFFSR_267 ( );
FILL FILL_4_DFFSR_267 ( );
FILL FILL_5_DFFSR_267 ( );
FILL FILL_6_DFFSR_267 ( );
FILL FILL_7_DFFSR_267 ( );
FILL FILL_8_DFFSR_267 ( );
FILL FILL_9_DFFSR_267 ( );
FILL FILL_10_DFFSR_267 ( );
FILL FILL_11_DFFSR_267 ( );
FILL FILL_12_DFFSR_267 ( );
FILL FILL_13_DFFSR_267 ( );
FILL FILL_14_DFFSR_267 ( );
FILL FILL_15_DFFSR_267 ( );
FILL FILL_16_DFFSR_267 ( );
FILL FILL_17_DFFSR_267 ( );
FILL FILL_18_DFFSR_267 ( );
FILL FILL_19_DFFSR_267 ( );
FILL FILL_20_DFFSR_267 ( );
FILL FILL_21_DFFSR_267 ( );
FILL FILL_22_DFFSR_267 ( );
FILL FILL_23_DFFSR_267 ( );
FILL FILL_24_DFFSR_267 ( );
FILL FILL_25_DFFSR_267 ( );
FILL FILL_26_DFFSR_267 ( );
FILL FILL_27_DFFSR_267 ( );
FILL FILL_28_DFFSR_267 ( );
FILL FILL_29_DFFSR_267 ( );
FILL FILL_30_DFFSR_267 ( );
FILL FILL_31_DFFSR_267 ( );
FILL FILL_32_DFFSR_267 ( );
FILL FILL_33_DFFSR_267 ( );
FILL FILL_34_DFFSR_267 ( );
FILL FILL_35_DFFSR_267 ( );
FILL FILL_36_DFFSR_267 ( );
FILL FILL_37_DFFSR_267 ( );
FILL FILL_38_DFFSR_267 ( );
FILL FILL_39_DFFSR_267 ( );
FILL FILL_40_DFFSR_267 ( );
FILL FILL_41_DFFSR_267 ( );
FILL FILL_42_DFFSR_267 ( );
FILL FILL_43_DFFSR_267 ( );
FILL FILL_44_DFFSR_267 ( );
FILL FILL_45_DFFSR_267 ( );
FILL FILL_46_DFFSR_267 ( );
FILL FILL_47_DFFSR_267 ( );
FILL FILL_48_DFFSR_267 ( );
FILL FILL_49_DFFSR_267 ( );
FILL FILL_50_DFFSR_267 ( );
FILL FILL_0_OAI21X1_101 ( );
FILL FILL_1_OAI21X1_101 ( );
FILL FILL_2_OAI21X1_101 ( );
FILL FILL_3_OAI21X1_101 ( );
FILL FILL_4_OAI21X1_101 ( );
FILL FILL_5_OAI21X1_101 ( );
FILL FILL_6_OAI21X1_101 ( );
FILL FILL_7_OAI21X1_101 ( );
FILL FILL_8_OAI21X1_101 ( );
FILL FILL_0_DFFSR_182 ( );
FILL FILL_1_DFFSR_182 ( );
FILL FILL_2_DFFSR_182 ( );
FILL FILL_3_DFFSR_182 ( );
FILL FILL_4_DFFSR_182 ( );
FILL FILL_5_DFFSR_182 ( );
FILL FILL_6_DFFSR_182 ( );
FILL FILL_7_DFFSR_182 ( );
FILL FILL_8_DFFSR_182 ( );
FILL FILL_9_DFFSR_182 ( );
FILL FILL_10_DFFSR_182 ( );
FILL FILL_11_DFFSR_182 ( );
FILL FILL_12_DFFSR_182 ( );
FILL FILL_13_DFFSR_182 ( );
FILL FILL_14_DFFSR_182 ( );
FILL FILL_15_DFFSR_182 ( );
FILL FILL_16_DFFSR_182 ( );
FILL FILL_17_DFFSR_182 ( );
FILL FILL_18_DFFSR_182 ( );
FILL FILL_19_DFFSR_182 ( );
FILL FILL_20_DFFSR_182 ( );
FILL FILL_21_DFFSR_182 ( );
FILL FILL_22_DFFSR_182 ( );
FILL FILL_23_DFFSR_182 ( );
FILL FILL_24_DFFSR_182 ( );
FILL FILL_25_DFFSR_182 ( );
FILL FILL_26_DFFSR_182 ( );
FILL FILL_27_DFFSR_182 ( );
FILL FILL_28_DFFSR_182 ( );
FILL FILL_29_DFFSR_182 ( );
FILL FILL_30_DFFSR_182 ( );
FILL FILL_31_DFFSR_182 ( );
FILL FILL_32_DFFSR_182 ( );
FILL FILL_33_DFFSR_182 ( );
FILL FILL_34_DFFSR_182 ( );
FILL FILL_35_DFFSR_182 ( );
FILL FILL_36_DFFSR_182 ( );
FILL FILL_37_DFFSR_182 ( );
FILL FILL_38_DFFSR_182 ( );
FILL FILL_39_DFFSR_182 ( );
FILL FILL_40_DFFSR_182 ( );
FILL FILL_41_DFFSR_182 ( );
FILL FILL_42_DFFSR_182 ( );
FILL FILL_43_DFFSR_182 ( );
FILL FILL_44_DFFSR_182 ( );
FILL FILL_45_DFFSR_182 ( );
FILL FILL_46_DFFSR_182 ( );
FILL FILL_47_DFFSR_182 ( );
FILL FILL_48_DFFSR_182 ( );
FILL FILL_49_DFFSR_182 ( );
FILL FILL_50_DFFSR_182 ( );
FILL FILL_51_DFFSR_182 ( );
FILL FILL_0_DFFSR_228 ( );
FILL FILL_1_DFFSR_228 ( );
FILL FILL_2_DFFSR_228 ( );
FILL FILL_3_DFFSR_228 ( );
FILL FILL_4_DFFSR_228 ( );
FILL FILL_5_DFFSR_228 ( );
FILL FILL_6_DFFSR_228 ( );
FILL FILL_7_DFFSR_228 ( );
FILL FILL_8_DFFSR_228 ( );
FILL FILL_9_DFFSR_228 ( );
FILL FILL_10_DFFSR_228 ( );
FILL FILL_11_DFFSR_228 ( );
FILL FILL_12_DFFSR_228 ( );
FILL FILL_13_DFFSR_228 ( );
FILL FILL_14_DFFSR_228 ( );
FILL FILL_15_DFFSR_228 ( );
FILL FILL_16_DFFSR_228 ( );
FILL FILL_17_DFFSR_228 ( );
FILL FILL_18_DFFSR_228 ( );
FILL FILL_19_DFFSR_228 ( );
FILL FILL_20_DFFSR_228 ( );
FILL FILL_21_DFFSR_228 ( );
FILL FILL_22_DFFSR_228 ( );
FILL FILL_23_DFFSR_228 ( );
FILL FILL_24_DFFSR_228 ( );
FILL FILL_25_DFFSR_228 ( );
FILL FILL_26_DFFSR_228 ( );
FILL FILL_27_DFFSR_228 ( );
FILL FILL_28_DFFSR_228 ( );
FILL FILL_29_DFFSR_228 ( );
FILL FILL_30_DFFSR_228 ( );
FILL FILL_31_DFFSR_228 ( );
FILL FILL_32_DFFSR_228 ( );
FILL FILL_33_DFFSR_228 ( );
FILL FILL_34_DFFSR_228 ( );
FILL FILL_35_DFFSR_228 ( );
FILL FILL_36_DFFSR_228 ( );
FILL FILL_37_DFFSR_228 ( );
FILL FILL_38_DFFSR_228 ( );
FILL FILL_39_DFFSR_228 ( );
FILL FILL_40_DFFSR_228 ( );
FILL FILL_41_DFFSR_228 ( );
FILL FILL_42_DFFSR_228 ( );
FILL FILL_43_DFFSR_228 ( );
FILL FILL_44_DFFSR_228 ( );
FILL FILL_45_DFFSR_228 ( );
FILL FILL_46_DFFSR_228 ( );
FILL FILL_47_DFFSR_228 ( );
FILL FILL_48_DFFSR_228 ( );
FILL FILL_49_DFFSR_228 ( );
FILL FILL_50_DFFSR_228 ( );
FILL FILL_0_AOI22X1_12 ( );
FILL FILL_1_AOI22X1_12 ( );
FILL FILL_2_AOI22X1_12 ( );
FILL FILL_3_AOI22X1_12 ( );
FILL FILL_4_AOI22X1_12 ( );
FILL FILL_5_AOI22X1_12 ( );
FILL FILL_6_AOI22X1_12 ( );
FILL FILL_7_AOI22X1_12 ( );
FILL FILL_8_AOI22X1_12 ( );
FILL FILL_9_AOI22X1_12 ( );
FILL FILL_10_AOI22X1_12 ( );
FILL FILL_11_AOI22X1_12 ( );
FILL FILL_0_BUFX2_68 ( );
FILL FILL_1_BUFX2_68 ( );
FILL FILL_2_BUFX2_68 ( );
FILL FILL_3_BUFX2_68 ( );
FILL FILL_4_BUFX2_68 ( );
FILL FILL_5_BUFX2_68 ( );
FILL FILL_6_BUFX2_68 ( );
FILL FILL_0_NAND3X1_93 ( );
FILL FILL_1_NAND3X1_93 ( );
FILL FILL_2_NAND3X1_93 ( );
FILL FILL_3_NAND3X1_93 ( );
FILL FILL_4_NAND3X1_93 ( );
FILL FILL_5_NAND3X1_93 ( );
FILL FILL_6_NAND3X1_93 ( );
FILL FILL_7_NAND3X1_93 ( );
FILL FILL_8_NAND3X1_93 ( );
FILL FILL_9_NAND3X1_93 ( );
FILL FILL_0_DFFSR_246 ( );
FILL FILL_1_DFFSR_246 ( );
FILL FILL_2_DFFSR_246 ( );
FILL FILL_3_DFFSR_246 ( );
FILL FILL_4_DFFSR_246 ( );
FILL FILL_5_DFFSR_246 ( );
FILL FILL_6_DFFSR_246 ( );
FILL FILL_7_DFFSR_246 ( );
FILL FILL_8_DFFSR_246 ( );
FILL FILL_9_DFFSR_246 ( );
FILL FILL_10_DFFSR_246 ( );
FILL FILL_11_DFFSR_246 ( );
FILL FILL_12_DFFSR_246 ( );
FILL FILL_13_DFFSR_246 ( );
FILL FILL_14_DFFSR_246 ( );
FILL FILL_15_DFFSR_246 ( );
FILL FILL_16_DFFSR_246 ( );
FILL FILL_17_DFFSR_246 ( );
FILL FILL_18_DFFSR_246 ( );
FILL FILL_19_DFFSR_246 ( );
FILL FILL_20_DFFSR_246 ( );
FILL FILL_21_DFFSR_246 ( );
FILL FILL_22_DFFSR_246 ( );
FILL FILL_23_DFFSR_246 ( );
FILL FILL_24_DFFSR_246 ( );
FILL FILL_25_DFFSR_246 ( );
FILL FILL_26_DFFSR_246 ( );
FILL FILL_27_DFFSR_246 ( );
FILL FILL_28_DFFSR_246 ( );
FILL FILL_29_DFFSR_246 ( );
FILL FILL_30_DFFSR_246 ( );
FILL FILL_31_DFFSR_246 ( );
FILL FILL_32_DFFSR_246 ( );
FILL FILL_33_DFFSR_246 ( );
FILL FILL_34_DFFSR_246 ( );
FILL FILL_35_DFFSR_246 ( );
FILL FILL_36_DFFSR_246 ( );
FILL FILL_37_DFFSR_246 ( );
FILL FILL_38_DFFSR_246 ( );
FILL FILL_39_DFFSR_246 ( );
FILL FILL_40_DFFSR_246 ( );
FILL FILL_41_DFFSR_246 ( );
FILL FILL_42_DFFSR_246 ( );
FILL FILL_43_DFFSR_246 ( );
FILL FILL_44_DFFSR_246 ( );
FILL FILL_45_DFFSR_246 ( );
FILL FILL_46_DFFSR_246 ( );
FILL FILL_47_DFFSR_246 ( );
FILL FILL_48_DFFSR_246 ( );
FILL FILL_49_DFFSR_246 ( );
FILL FILL_50_DFFSR_246 ( );
FILL FILL_0_OAI21X1_11 ( );
FILL FILL_1_OAI21X1_11 ( );
FILL FILL_2_OAI21X1_11 ( );
FILL FILL_3_OAI21X1_11 ( );
FILL FILL_4_OAI21X1_11 ( );
FILL FILL_5_OAI21X1_11 ( );
FILL FILL_6_OAI21X1_11 ( );
FILL FILL_7_OAI21X1_11 ( );
FILL FILL_8_OAI21X1_11 ( );
FILL FILL_0_NAND3X1_114 ( );
FILL FILL_1_NAND3X1_114 ( );
FILL FILL_2_NAND3X1_114 ( );
FILL FILL_3_NAND3X1_114 ( );
FILL FILL_4_NAND3X1_114 ( );
FILL FILL_5_NAND3X1_114 ( );
FILL FILL_6_NAND3X1_114 ( );
FILL FILL_7_NAND3X1_114 ( );
FILL FILL_8_NAND3X1_114 ( );
FILL FILL_0_DFFSR_199 ( );
FILL FILL_1_DFFSR_199 ( );
FILL FILL_2_DFFSR_199 ( );
FILL FILL_3_DFFSR_199 ( );
FILL FILL_4_DFFSR_199 ( );
FILL FILL_5_DFFSR_199 ( );
FILL FILL_6_DFFSR_199 ( );
FILL FILL_7_DFFSR_199 ( );
FILL FILL_8_DFFSR_199 ( );
FILL FILL_9_DFFSR_199 ( );
FILL FILL_10_DFFSR_199 ( );
FILL FILL_11_DFFSR_199 ( );
FILL FILL_12_DFFSR_199 ( );
FILL FILL_13_DFFSR_199 ( );
FILL FILL_14_DFFSR_199 ( );
FILL FILL_15_DFFSR_199 ( );
FILL FILL_16_DFFSR_199 ( );
FILL FILL_17_DFFSR_199 ( );
FILL FILL_18_DFFSR_199 ( );
FILL FILL_19_DFFSR_199 ( );
FILL FILL_20_DFFSR_199 ( );
FILL FILL_21_DFFSR_199 ( );
FILL FILL_22_DFFSR_199 ( );
FILL FILL_23_DFFSR_199 ( );
FILL FILL_24_DFFSR_199 ( );
FILL FILL_25_DFFSR_199 ( );
FILL FILL_26_DFFSR_199 ( );
FILL FILL_27_DFFSR_199 ( );
FILL FILL_28_DFFSR_199 ( );
FILL FILL_29_DFFSR_199 ( );
FILL FILL_30_DFFSR_199 ( );
FILL FILL_31_DFFSR_199 ( );
FILL FILL_32_DFFSR_199 ( );
FILL FILL_33_DFFSR_199 ( );
FILL FILL_34_DFFSR_199 ( );
FILL FILL_35_DFFSR_199 ( );
FILL FILL_36_DFFSR_199 ( );
FILL FILL_37_DFFSR_199 ( );
FILL FILL_38_DFFSR_199 ( );
FILL FILL_39_DFFSR_199 ( );
FILL FILL_40_DFFSR_199 ( );
FILL FILL_41_DFFSR_199 ( );
FILL FILL_42_DFFSR_199 ( );
FILL FILL_43_DFFSR_199 ( );
FILL FILL_44_DFFSR_199 ( );
FILL FILL_45_DFFSR_199 ( );
FILL FILL_46_DFFSR_199 ( );
FILL FILL_47_DFFSR_199 ( );
FILL FILL_48_DFFSR_199 ( );
FILL FILL_49_DFFSR_199 ( );
FILL FILL_50_DFFSR_199 ( );
FILL FILL_51_DFFSR_199 ( );
FILL FILL_0_DFFSR_173 ( );
FILL FILL_1_DFFSR_173 ( );
FILL FILL_2_DFFSR_173 ( );
FILL FILL_3_DFFSR_173 ( );
FILL FILL_4_DFFSR_173 ( );
FILL FILL_5_DFFSR_173 ( );
FILL FILL_6_DFFSR_173 ( );
FILL FILL_7_DFFSR_173 ( );
FILL FILL_8_DFFSR_173 ( );
FILL FILL_9_DFFSR_173 ( );
FILL FILL_10_DFFSR_173 ( );
FILL FILL_11_DFFSR_173 ( );
FILL FILL_12_DFFSR_173 ( );
FILL FILL_13_DFFSR_173 ( );
FILL FILL_14_DFFSR_173 ( );
FILL FILL_15_DFFSR_173 ( );
FILL FILL_16_DFFSR_173 ( );
FILL FILL_17_DFFSR_173 ( );
FILL FILL_18_DFFSR_173 ( );
FILL FILL_19_DFFSR_173 ( );
FILL FILL_20_DFFSR_173 ( );
FILL FILL_21_DFFSR_173 ( );
FILL FILL_22_DFFSR_173 ( );
FILL FILL_23_DFFSR_173 ( );
FILL FILL_24_DFFSR_173 ( );
FILL FILL_25_DFFSR_173 ( );
FILL FILL_26_DFFSR_173 ( );
FILL FILL_27_DFFSR_173 ( );
FILL FILL_28_DFFSR_173 ( );
FILL FILL_29_DFFSR_173 ( );
FILL FILL_30_DFFSR_173 ( );
FILL FILL_31_DFFSR_173 ( );
FILL FILL_32_DFFSR_173 ( );
FILL FILL_33_DFFSR_173 ( );
FILL FILL_34_DFFSR_173 ( );
FILL FILL_35_DFFSR_173 ( );
FILL FILL_36_DFFSR_173 ( );
FILL FILL_37_DFFSR_173 ( );
FILL FILL_38_DFFSR_173 ( );
FILL FILL_39_DFFSR_173 ( );
FILL FILL_40_DFFSR_173 ( );
FILL FILL_41_DFFSR_173 ( );
FILL FILL_42_DFFSR_173 ( );
FILL FILL_43_DFFSR_173 ( );
FILL FILL_44_DFFSR_173 ( );
FILL FILL_45_DFFSR_173 ( );
FILL FILL_46_DFFSR_173 ( );
FILL FILL_47_DFFSR_173 ( );
FILL FILL_48_DFFSR_173 ( );
FILL FILL_49_DFFSR_173 ( );
FILL FILL_50_DFFSR_173 ( );
FILL FILL_51_DFFSR_173 ( );
FILL FILL_0_OAI21X1_51 ( );
FILL FILL_1_OAI21X1_51 ( );
FILL FILL_2_OAI21X1_51 ( );
FILL FILL_3_OAI21X1_51 ( );
FILL FILL_4_OAI21X1_51 ( );
FILL FILL_5_OAI21X1_51 ( );
FILL FILL_6_OAI21X1_51 ( );
FILL FILL_7_OAI21X1_51 ( );
FILL FILL_8_OAI21X1_51 ( );
FILL FILL_0_AOI21X1_32 ( );
FILL FILL_1_AOI21X1_32 ( );
FILL FILL_2_AOI21X1_32 ( );
FILL FILL_3_AOI21X1_32 ( );
FILL FILL_4_AOI21X1_32 ( );
FILL FILL_5_AOI21X1_32 ( );
FILL FILL_6_AOI21X1_32 ( );
FILL FILL_7_AOI21X1_32 ( );
FILL FILL_8_AOI21X1_32 ( );
FILL FILL_9_AOI21X1_32 ( );
FILL FILL_0_AOI21X1_29 ( );
FILL FILL_1_AOI21X1_29 ( );
FILL FILL_2_AOI21X1_29 ( );
FILL FILL_3_AOI21X1_29 ( );
FILL FILL_4_AOI21X1_29 ( );
FILL FILL_5_AOI21X1_29 ( );
FILL FILL_6_AOI21X1_29 ( );
FILL FILL_7_AOI21X1_29 ( );
FILL FILL_8_AOI21X1_29 ( );
FILL FILL_0_OAI21X1_59 ( );
FILL FILL_1_OAI21X1_59 ( );
FILL FILL_2_OAI21X1_59 ( );
FILL FILL_3_OAI21X1_59 ( );
FILL FILL_4_OAI21X1_59 ( );
FILL FILL_5_OAI21X1_59 ( );
FILL FILL_6_OAI21X1_59 ( );
FILL FILL_7_OAI21X1_59 ( );
FILL FILL_8_OAI21X1_59 ( );
FILL FILL_0_AOI21X1_26 ( );
FILL FILL_1_AOI21X1_26 ( );
FILL FILL_2_AOI21X1_26 ( );
FILL FILL_3_AOI21X1_26 ( );
FILL FILL_4_AOI21X1_26 ( );
FILL FILL_5_AOI21X1_26 ( );
FILL FILL_6_AOI21X1_26 ( );
FILL FILL_7_AOI21X1_26 ( );
FILL FILL_8_AOI21X1_26 ( );
FILL FILL_0_AOI21X1_25 ( );
FILL FILL_1_AOI21X1_25 ( );
FILL FILL_2_AOI21X1_25 ( );
FILL FILL_3_AOI21X1_25 ( );
FILL FILL_4_AOI21X1_25 ( );
FILL FILL_5_AOI21X1_25 ( );
FILL FILL_6_AOI21X1_25 ( );
FILL FILL_7_AOI21X1_25 ( );
FILL FILL_8_AOI21X1_25 ( );
FILL FILL_0_NAND2X1_59 ( );
FILL FILL_1_NAND2X1_59 ( );
FILL FILL_2_NAND2X1_59 ( );
FILL FILL_3_NAND2X1_59 ( );
FILL FILL_4_NAND2X1_59 ( );
FILL FILL_5_NAND2X1_59 ( );
FILL FILL_6_NAND2X1_59 ( );
FILL FILL_0_NAND3X1_194 ( );
FILL FILL_1_NAND3X1_194 ( );
FILL FILL_2_NAND3X1_194 ( );
FILL FILL_3_NAND3X1_194 ( );
FILL FILL_4_NAND3X1_194 ( );
FILL FILL_5_NAND3X1_194 ( );
FILL FILL_6_NAND3X1_194 ( );
FILL FILL_7_NAND3X1_194 ( );
FILL FILL_8_NAND3X1_194 ( );
FILL FILL_9_NAND3X1_194 ( );
FILL FILL_0_AOI21X1_19 ( );
FILL FILL_1_AOI21X1_19 ( );
FILL FILL_2_AOI21X1_19 ( );
FILL FILL_3_AOI21X1_19 ( );
FILL FILL_4_AOI21X1_19 ( );
FILL FILL_5_AOI21X1_19 ( );
FILL FILL_6_AOI21X1_19 ( );
FILL FILL_7_AOI21X1_19 ( );
FILL FILL_8_AOI21X1_19 ( );
FILL FILL_0_OAI21X1_55 ( );
FILL FILL_1_OAI21X1_55 ( );
FILL FILL_2_OAI21X1_55 ( );
FILL FILL_3_OAI21X1_55 ( );
FILL FILL_4_OAI21X1_55 ( );
FILL FILL_5_OAI21X1_55 ( );
FILL FILL_6_OAI21X1_55 ( );
FILL FILL_7_OAI21X1_55 ( );
FILL FILL_8_OAI21X1_55 ( );
FILL FILL_0_OAI21X1_44 ( );
FILL FILL_1_OAI21X1_44 ( );
FILL FILL_2_OAI21X1_44 ( );
FILL FILL_3_OAI21X1_44 ( );
FILL FILL_4_OAI21X1_44 ( );
FILL FILL_5_OAI21X1_44 ( );
FILL FILL_6_OAI21X1_44 ( );
FILL FILL_7_OAI21X1_44 ( );
FILL FILL_8_OAI21X1_44 ( );
FILL FILL_9_OAI21X1_44 ( );
FILL FILL_0_OAI21X1_45 ( );
FILL FILL_1_OAI21X1_45 ( );
FILL FILL_2_OAI21X1_45 ( );
FILL FILL_3_OAI21X1_45 ( );
FILL FILL_4_OAI21X1_45 ( );
FILL FILL_5_OAI21X1_45 ( );
FILL FILL_6_OAI21X1_45 ( );
FILL FILL_7_OAI21X1_45 ( );
FILL FILL_8_OAI21X1_45 ( );
FILL FILL_0_NOR2X1_74 ( );
FILL FILL_1_NOR2X1_74 ( );
FILL FILL_2_NOR2X1_74 ( );
FILL FILL_3_NOR2X1_74 ( );
FILL FILL_4_NOR2X1_74 ( );
FILL FILL_5_NOR2X1_74 ( );
FILL FILL_6_NOR2X1_74 ( );
FILL FILL_0_NAND2X1_165 ( );
FILL FILL_1_NAND2X1_165 ( );
FILL FILL_2_NAND2X1_165 ( );
FILL FILL_3_NAND2X1_165 ( );
FILL FILL_4_NAND2X1_165 ( );
FILL FILL_5_NAND2X1_165 ( );
FILL FILL_6_NAND2X1_165 ( );
FILL FILL_0_INVX1_120 ( );
FILL FILL_1_INVX1_120 ( );
FILL FILL_2_INVX1_120 ( );
FILL FILL_3_INVX1_120 ( );
FILL FILL_4_INVX1_120 ( );
FILL FILL_0_AOI21X1_2 ( );
FILL FILL_1_AOI21X1_2 ( );
FILL FILL_2_AOI21X1_2 ( );
FILL FILL_3_AOI21X1_2 ( );
FILL FILL_4_AOI21X1_2 ( );
FILL FILL_5_AOI21X1_2 ( );
FILL FILL_6_AOI21X1_2 ( );
FILL FILL_7_AOI21X1_2 ( );
FILL FILL_8_AOI21X1_2 ( );
FILL FILL_0_DFFSR_273 ( );
FILL FILL_1_DFFSR_273 ( );
FILL FILL_2_DFFSR_273 ( );
FILL FILL_3_DFFSR_273 ( );
FILL FILL_4_DFFSR_273 ( );
FILL FILL_5_DFFSR_273 ( );
FILL FILL_6_DFFSR_273 ( );
FILL FILL_7_DFFSR_273 ( );
FILL FILL_8_DFFSR_273 ( );
FILL FILL_9_DFFSR_273 ( );
FILL FILL_10_DFFSR_273 ( );
FILL FILL_11_DFFSR_273 ( );
FILL FILL_12_DFFSR_273 ( );
FILL FILL_13_DFFSR_273 ( );
FILL FILL_14_DFFSR_273 ( );
FILL FILL_15_DFFSR_273 ( );
FILL FILL_16_DFFSR_273 ( );
FILL FILL_17_DFFSR_273 ( );
FILL FILL_18_DFFSR_273 ( );
FILL FILL_19_DFFSR_273 ( );
FILL FILL_20_DFFSR_273 ( );
FILL FILL_21_DFFSR_273 ( );
FILL FILL_22_DFFSR_273 ( );
FILL FILL_23_DFFSR_273 ( );
FILL FILL_24_DFFSR_273 ( );
FILL FILL_25_DFFSR_273 ( );
FILL FILL_26_DFFSR_273 ( );
FILL FILL_27_DFFSR_273 ( );
FILL FILL_28_DFFSR_273 ( );
FILL FILL_29_DFFSR_273 ( );
FILL FILL_30_DFFSR_273 ( );
FILL FILL_31_DFFSR_273 ( );
FILL FILL_32_DFFSR_273 ( );
FILL FILL_33_DFFSR_273 ( );
FILL FILL_34_DFFSR_273 ( );
FILL FILL_35_DFFSR_273 ( );
FILL FILL_36_DFFSR_273 ( );
FILL FILL_37_DFFSR_273 ( );
FILL FILL_38_DFFSR_273 ( );
FILL FILL_39_DFFSR_273 ( );
FILL FILL_40_DFFSR_273 ( );
FILL FILL_41_DFFSR_273 ( );
FILL FILL_42_DFFSR_273 ( );
FILL FILL_43_DFFSR_273 ( );
FILL FILL_44_DFFSR_273 ( );
FILL FILL_45_DFFSR_273 ( );
FILL FILL_46_DFFSR_273 ( );
FILL FILL_47_DFFSR_273 ( );
FILL FILL_48_DFFSR_273 ( );
FILL FILL_49_DFFSR_273 ( );
FILL FILL_50_DFFSR_273 ( );
FILL FILL_0_DFFSR_135 ( );
FILL FILL_1_DFFSR_135 ( );
FILL FILL_2_DFFSR_135 ( );
FILL FILL_3_DFFSR_135 ( );
FILL FILL_4_DFFSR_135 ( );
FILL FILL_5_DFFSR_135 ( );
FILL FILL_6_DFFSR_135 ( );
FILL FILL_7_DFFSR_135 ( );
FILL FILL_8_DFFSR_135 ( );
FILL FILL_9_DFFSR_135 ( );
FILL FILL_10_DFFSR_135 ( );
FILL FILL_11_DFFSR_135 ( );
FILL FILL_12_DFFSR_135 ( );
FILL FILL_13_DFFSR_135 ( );
FILL FILL_14_DFFSR_135 ( );
FILL FILL_15_DFFSR_135 ( );
FILL FILL_16_DFFSR_135 ( );
FILL FILL_17_DFFSR_135 ( );
FILL FILL_18_DFFSR_135 ( );
FILL FILL_19_DFFSR_135 ( );
FILL FILL_20_DFFSR_135 ( );
FILL FILL_21_DFFSR_135 ( );
FILL FILL_22_DFFSR_135 ( );
FILL FILL_23_DFFSR_135 ( );
FILL FILL_24_DFFSR_135 ( );
FILL FILL_25_DFFSR_135 ( );
FILL FILL_26_DFFSR_135 ( );
FILL FILL_27_DFFSR_135 ( );
FILL FILL_28_DFFSR_135 ( );
FILL FILL_29_DFFSR_135 ( );
FILL FILL_30_DFFSR_135 ( );
FILL FILL_31_DFFSR_135 ( );
FILL FILL_32_DFFSR_135 ( );
FILL FILL_33_DFFSR_135 ( );
FILL FILL_34_DFFSR_135 ( );
FILL FILL_35_DFFSR_135 ( );
FILL FILL_36_DFFSR_135 ( );
FILL FILL_37_DFFSR_135 ( );
FILL FILL_38_DFFSR_135 ( );
FILL FILL_39_DFFSR_135 ( );
FILL FILL_40_DFFSR_135 ( );
FILL FILL_41_DFFSR_135 ( );
FILL FILL_42_DFFSR_135 ( );
FILL FILL_43_DFFSR_135 ( );
FILL FILL_44_DFFSR_135 ( );
FILL FILL_45_DFFSR_135 ( );
FILL FILL_46_DFFSR_135 ( );
FILL FILL_47_DFFSR_135 ( );
FILL FILL_48_DFFSR_135 ( );
FILL FILL_49_DFFSR_135 ( );
FILL FILL_50_DFFSR_135 ( );
FILL FILL_0_DFFSR_140 ( );
FILL FILL_1_DFFSR_140 ( );
FILL FILL_2_DFFSR_140 ( );
FILL FILL_3_DFFSR_140 ( );
FILL FILL_4_DFFSR_140 ( );
FILL FILL_5_DFFSR_140 ( );
FILL FILL_6_DFFSR_140 ( );
FILL FILL_7_DFFSR_140 ( );
FILL FILL_8_DFFSR_140 ( );
FILL FILL_9_DFFSR_140 ( );
FILL FILL_10_DFFSR_140 ( );
FILL FILL_11_DFFSR_140 ( );
FILL FILL_12_DFFSR_140 ( );
FILL FILL_13_DFFSR_140 ( );
FILL FILL_14_DFFSR_140 ( );
FILL FILL_15_DFFSR_140 ( );
FILL FILL_16_DFFSR_140 ( );
FILL FILL_17_DFFSR_140 ( );
FILL FILL_18_DFFSR_140 ( );
FILL FILL_19_DFFSR_140 ( );
FILL FILL_20_DFFSR_140 ( );
FILL FILL_21_DFFSR_140 ( );
FILL FILL_22_DFFSR_140 ( );
FILL FILL_23_DFFSR_140 ( );
FILL FILL_24_DFFSR_140 ( );
FILL FILL_25_DFFSR_140 ( );
FILL FILL_26_DFFSR_140 ( );
FILL FILL_27_DFFSR_140 ( );
FILL FILL_28_DFFSR_140 ( );
FILL FILL_29_DFFSR_140 ( );
FILL FILL_30_DFFSR_140 ( );
FILL FILL_31_DFFSR_140 ( );
FILL FILL_32_DFFSR_140 ( );
FILL FILL_33_DFFSR_140 ( );
FILL FILL_34_DFFSR_140 ( );
FILL FILL_35_DFFSR_140 ( );
FILL FILL_36_DFFSR_140 ( );
FILL FILL_37_DFFSR_140 ( );
FILL FILL_38_DFFSR_140 ( );
FILL FILL_39_DFFSR_140 ( );
FILL FILL_40_DFFSR_140 ( );
FILL FILL_41_DFFSR_140 ( );
FILL FILL_42_DFFSR_140 ( );
FILL FILL_43_DFFSR_140 ( );
FILL FILL_44_DFFSR_140 ( );
FILL FILL_45_DFFSR_140 ( );
FILL FILL_46_DFFSR_140 ( );
FILL FILL_47_DFFSR_140 ( );
FILL FILL_48_DFFSR_140 ( );
FILL FILL_49_DFFSR_140 ( );
FILL FILL_50_DFFSR_140 ( );
FILL FILL_51_DFFSR_140 ( );
FILL FILL_0_NAND3X1_94 ( );
FILL FILL_1_NAND3X1_94 ( );
FILL FILL_2_NAND3X1_94 ( );
FILL FILL_3_NAND3X1_94 ( );
FILL FILL_4_NAND3X1_94 ( );
FILL FILL_5_NAND3X1_94 ( );
FILL FILL_6_NAND3X1_94 ( );
FILL FILL_7_NAND3X1_94 ( );
FILL FILL_8_NAND3X1_94 ( );
FILL FILL_0_NAND3X1_95 ( );
FILL FILL_1_NAND3X1_95 ( );
FILL FILL_2_NAND3X1_95 ( );
FILL FILL_3_NAND3X1_95 ( );
FILL FILL_4_NAND3X1_95 ( );
FILL FILL_5_NAND3X1_95 ( );
FILL FILL_6_NAND3X1_95 ( );
FILL FILL_7_NAND3X1_95 ( );
FILL FILL_8_NAND3X1_95 ( );
FILL FILL_0_BUFX2_27 ( );
FILL FILL_1_BUFX2_27 ( );
FILL FILL_2_BUFX2_27 ( );
FILL FILL_3_BUFX2_27 ( );
FILL FILL_4_BUFX2_27 ( );
FILL FILL_5_BUFX2_27 ( );
FILL FILL_6_BUFX2_27 ( );
FILL FILL_0_NAND3X1_65 ( );
FILL FILL_1_NAND3X1_65 ( );
FILL FILL_2_NAND3X1_65 ( );
FILL FILL_3_NAND3X1_65 ( );
FILL FILL_4_NAND3X1_65 ( );
FILL FILL_5_NAND3X1_65 ( );
FILL FILL_6_NAND3X1_65 ( );
FILL FILL_7_NAND3X1_65 ( );
FILL FILL_8_NAND3X1_65 ( );
FILL FILL_9_NAND3X1_65 ( );
FILL FILL_0_NAND2X1_47 ( );
FILL FILL_1_NAND2X1_47 ( );
FILL FILL_2_NAND2X1_47 ( );
FILL FILL_3_NAND2X1_47 ( );
FILL FILL_4_NAND2X1_47 ( );
FILL FILL_5_NAND2X1_47 ( );
FILL FILL_6_NAND2X1_47 ( );
FILL FILL_0_OAI21X1_14 ( );
FILL FILL_1_OAI21X1_14 ( );
FILL FILL_2_OAI21X1_14 ( );
FILL FILL_3_OAI21X1_14 ( );
FILL FILL_4_OAI21X1_14 ( );
FILL FILL_5_OAI21X1_14 ( );
FILL FILL_6_OAI21X1_14 ( );
FILL FILL_7_OAI21X1_14 ( );
FILL FILL_8_OAI21X1_14 ( );
FILL FILL_0_DFFSR_159 ( );
FILL FILL_1_DFFSR_159 ( );
FILL FILL_2_DFFSR_159 ( );
FILL FILL_3_DFFSR_159 ( );
FILL FILL_4_DFFSR_159 ( );
FILL FILL_5_DFFSR_159 ( );
FILL FILL_6_DFFSR_159 ( );
FILL FILL_7_DFFSR_159 ( );
FILL FILL_8_DFFSR_159 ( );
FILL FILL_9_DFFSR_159 ( );
FILL FILL_10_DFFSR_159 ( );
FILL FILL_11_DFFSR_159 ( );
FILL FILL_12_DFFSR_159 ( );
FILL FILL_13_DFFSR_159 ( );
FILL FILL_14_DFFSR_159 ( );
FILL FILL_15_DFFSR_159 ( );
FILL FILL_16_DFFSR_159 ( );
FILL FILL_17_DFFSR_159 ( );
FILL FILL_18_DFFSR_159 ( );
FILL FILL_19_DFFSR_159 ( );
FILL FILL_20_DFFSR_159 ( );
FILL FILL_21_DFFSR_159 ( );
FILL FILL_22_DFFSR_159 ( );
FILL FILL_23_DFFSR_159 ( );
FILL FILL_24_DFFSR_159 ( );
FILL FILL_25_DFFSR_159 ( );
FILL FILL_26_DFFSR_159 ( );
FILL FILL_27_DFFSR_159 ( );
FILL FILL_28_DFFSR_159 ( );
FILL FILL_29_DFFSR_159 ( );
FILL FILL_30_DFFSR_159 ( );
FILL FILL_31_DFFSR_159 ( );
FILL FILL_32_DFFSR_159 ( );
FILL FILL_33_DFFSR_159 ( );
FILL FILL_34_DFFSR_159 ( );
FILL FILL_35_DFFSR_159 ( );
FILL FILL_36_DFFSR_159 ( );
FILL FILL_37_DFFSR_159 ( );
FILL FILL_38_DFFSR_159 ( );
FILL FILL_39_DFFSR_159 ( );
FILL FILL_40_DFFSR_159 ( );
FILL FILL_41_DFFSR_159 ( );
FILL FILL_42_DFFSR_159 ( );
FILL FILL_43_DFFSR_159 ( );
FILL FILL_44_DFFSR_159 ( );
FILL FILL_45_DFFSR_159 ( );
FILL FILL_46_DFFSR_159 ( );
FILL FILL_47_DFFSR_159 ( );
FILL FILL_48_DFFSR_159 ( );
FILL FILL_49_DFFSR_159 ( );
FILL FILL_50_DFFSR_159 ( );
FILL FILL_0_NAND3X1_117 ( );
FILL FILL_1_NAND3X1_117 ( );
FILL FILL_2_NAND3X1_117 ( );
FILL FILL_3_NAND3X1_117 ( );
FILL FILL_4_NAND3X1_117 ( );
FILL FILL_5_NAND3X1_117 ( );
FILL FILL_6_NAND3X1_117 ( );
FILL FILL_7_NAND3X1_117 ( );
FILL FILL_8_NAND3X1_117 ( );
FILL FILL_9_NAND3X1_117 ( );
FILL FILL_0_OAI22X1_43 ( );
FILL FILL_1_OAI22X1_43 ( );
FILL FILL_2_OAI22X1_43 ( );
FILL FILL_3_OAI22X1_43 ( );
FILL FILL_4_OAI22X1_43 ( );
FILL FILL_5_OAI22X1_43 ( );
FILL FILL_6_OAI22X1_43 ( );
FILL FILL_7_OAI22X1_43 ( );
FILL FILL_8_OAI22X1_43 ( );
FILL FILL_9_OAI22X1_43 ( );
FILL FILL_10_OAI22X1_43 ( );
FILL FILL_11_OAI22X1_43 ( );
FILL FILL_0_NAND3X1_113 ( );
FILL FILL_1_NAND3X1_113 ( );
FILL FILL_2_NAND3X1_113 ( );
FILL FILL_3_NAND3X1_113 ( );
FILL FILL_4_NAND3X1_113 ( );
FILL FILL_5_NAND3X1_113 ( );
FILL FILL_6_NAND3X1_113 ( );
FILL FILL_7_NAND3X1_113 ( );
FILL FILL_8_NAND3X1_113 ( );
FILL FILL_0_DFFSR_208 ( );
FILL FILL_1_DFFSR_208 ( );
FILL FILL_2_DFFSR_208 ( );
FILL FILL_3_DFFSR_208 ( );
FILL FILL_4_DFFSR_208 ( );
FILL FILL_5_DFFSR_208 ( );
FILL FILL_6_DFFSR_208 ( );
FILL FILL_7_DFFSR_208 ( );
FILL FILL_8_DFFSR_208 ( );
FILL FILL_9_DFFSR_208 ( );
FILL FILL_10_DFFSR_208 ( );
FILL FILL_11_DFFSR_208 ( );
FILL FILL_12_DFFSR_208 ( );
FILL FILL_13_DFFSR_208 ( );
FILL FILL_14_DFFSR_208 ( );
FILL FILL_15_DFFSR_208 ( );
FILL FILL_16_DFFSR_208 ( );
FILL FILL_17_DFFSR_208 ( );
FILL FILL_18_DFFSR_208 ( );
FILL FILL_19_DFFSR_208 ( );
FILL FILL_20_DFFSR_208 ( );
FILL FILL_21_DFFSR_208 ( );
FILL FILL_22_DFFSR_208 ( );
FILL FILL_23_DFFSR_208 ( );
FILL FILL_24_DFFSR_208 ( );
FILL FILL_25_DFFSR_208 ( );
FILL FILL_26_DFFSR_208 ( );
FILL FILL_27_DFFSR_208 ( );
FILL FILL_28_DFFSR_208 ( );
FILL FILL_29_DFFSR_208 ( );
FILL FILL_30_DFFSR_208 ( );
FILL FILL_31_DFFSR_208 ( );
FILL FILL_32_DFFSR_208 ( );
FILL FILL_33_DFFSR_208 ( );
FILL FILL_34_DFFSR_208 ( );
FILL FILL_35_DFFSR_208 ( );
FILL FILL_36_DFFSR_208 ( );
FILL FILL_37_DFFSR_208 ( );
FILL FILL_38_DFFSR_208 ( );
FILL FILL_39_DFFSR_208 ( );
FILL FILL_40_DFFSR_208 ( );
FILL FILL_41_DFFSR_208 ( );
FILL FILL_42_DFFSR_208 ( );
FILL FILL_43_DFFSR_208 ( );
FILL FILL_44_DFFSR_208 ( );
FILL FILL_45_DFFSR_208 ( );
FILL FILL_46_DFFSR_208 ( );
FILL FILL_47_DFFSR_208 ( );
FILL FILL_48_DFFSR_208 ( );
FILL FILL_49_DFFSR_208 ( );
FILL FILL_50_DFFSR_208 ( );
FILL FILL_51_DFFSR_208 ( );
FILL FILL_0_AOI21X1_22 ( );
FILL FILL_1_AOI21X1_22 ( );
FILL FILL_2_AOI21X1_22 ( );
FILL FILL_3_AOI21X1_22 ( );
FILL FILL_4_AOI21X1_22 ( );
FILL FILL_5_AOI21X1_22 ( );
FILL FILL_6_AOI21X1_22 ( );
FILL FILL_7_AOI21X1_22 ( );
FILL FILL_8_AOI21X1_22 ( );
FILL FILL_0_NAND3X1_198 ( );
FILL FILL_1_NAND3X1_198 ( );
FILL FILL_2_NAND3X1_198 ( );
FILL FILL_3_NAND3X1_198 ( );
FILL FILL_4_NAND3X1_198 ( );
FILL FILL_5_NAND3X1_198 ( );
FILL FILL_6_NAND3X1_198 ( );
FILL FILL_7_NAND3X1_198 ( );
FILL FILL_8_NAND3X1_198 ( );
FILL FILL_9_NAND3X1_198 ( );
FILL FILL_0_NAND3X1_215 ( );
FILL FILL_1_NAND3X1_215 ( );
FILL FILL_2_NAND3X1_215 ( );
FILL FILL_3_NAND3X1_215 ( );
FILL FILL_4_NAND3X1_215 ( );
FILL FILL_5_NAND3X1_215 ( );
FILL FILL_6_NAND3X1_215 ( );
FILL FILL_7_NAND3X1_215 ( );
FILL FILL_8_NAND3X1_215 ( );
FILL FILL_0_NAND3X1_219 ( );
FILL FILL_1_NAND3X1_219 ( );
FILL FILL_2_NAND3X1_219 ( );
FILL FILL_3_NAND3X1_219 ( );
FILL FILL_4_NAND3X1_219 ( );
FILL FILL_5_NAND3X1_219 ( );
FILL FILL_6_NAND3X1_219 ( );
FILL FILL_7_NAND3X1_219 ( );
FILL FILL_8_NAND3X1_219 ( );
FILL FILL_0_NAND2X1_137 ( );
FILL FILL_1_NAND2X1_137 ( );
FILL FILL_2_NAND2X1_137 ( );
FILL FILL_3_NAND2X1_137 ( );
FILL FILL_4_NAND2X1_137 ( );
FILL FILL_5_NAND2X1_137 ( );
FILL FILL_6_NAND2X1_137 ( );
FILL FILL_0_DFFPOSX1_14 ( );
FILL FILL_1_DFFPOSX1_14 ( );
FILL FILL_2_DFFPOSX1_14 ( );
FILL FILL_3_DFFPOSX1_14 ( );
FILL FILL_4_DFFPOSX1_14 ( );
FILL FILL_5_DFFPOSX1_14 ( );
FILL FILL_6_DFFPOSX1_14 ( );
FILL FILL_7_DFFPOSX1_14 ( );
FILL FILL_8_DFFPOSX1_14 ( );
FILL FILL_9_DFFPOSX1_14 ( );
FILL FILL_10_DFFPOSX1_14 ( );
FILL FILL_11_DFFPOSX1_14 ( );
FILL FILL_12_DFFPOSX1_14 ( );
FILL FILL_13_DFFPOSX1_14 ( );
FILL FILL_14_DFFPOSX1_14 ( );
FILL FILL_15_DFFPOSX1_14 ( );
FILL FILL_16_DFFPOSX1_14 ( );
FILL FILL_17_DFFPOSX1_14 ( );
FILL FILL_18_DFFPOSX1_14 ( );
FILL FILL_19_DFFPOSX1_14 ( );
FILL FILL_20_DFFPOSX1_14 ( );
FILL FILL_21_DFFPOSX1_14 ( );
FILL FILL_22_DFFPOSX1_14 ( );
FILL FILL_23_DFFPOSX1_14 ( );
FILL FILL_24_DFFPOSX1_14 ( );
FILL FILL_25_DFFPOSX1_14 ( );
FILL FILL_26_DFFPOSX1_14 ( );
FILL FILL_27_DFFPOSX1_14 ( );
FILL FILL_0_INVX1_142 ( );
FILL FILL_1_INVX1_142 ( );
FILL FILL_2_INVX1_142 ( );
FILL FILL_3_INVX1_142 ( );
FILL FILL_4_INVX1_142 ( );
FILL FILL_0_OAI21X1_25 ( );
FILL FILL_1_OAI21X1_25 ( );
FILL FILL_2_OAI21X1_25 ( );
FILL FILL_3_OAI21X1_25 ( );
FILL FILL_4_OAI21X1_25 ( );
FILL FILL_5_OAI21X1_25 ( );
FILL FILL_6_OAI21X1_25 ( );
FILL FILL_7_OAI21X1_25 ( );
FILL FILL_8_OAI21X1_25 ( );
FILL FILL_0_INVX1_156 ( );
FILL FILL_1_INVX1_156 ( );
FILL FILL_2_INVX1_156 ( );
FILL FILL_3_INVX1_156 ( );
FILL FILL_4_INVX1_156 ( );
FILL FILL_0_AOI21X1_23 ( );
FILL FILL_1_AOI21X1_23 ( );
FILL FILL_2_AOI21X1_23 ( );
FILL FILL_3_AOI21X1_23 ( );
FILL FILL_4_AOI21X1_23 ( );
FILL FILL_5_AOI21X1_23 ( );
FILL FILL_6_AOI21X1_23 ( );
FILL FILL_7_AOI21X1_23 ( );
FILL FILL_8_AOI21X1_23 ( );
FILL FILL_9_AOI21X1_23 ( );
FILL FILL_0_DFFPOSX1_4 ( );
FILL FILL_1_DFFPOSX1_4 ( );
FILL FILL_2_DFFPOSX1_4 ( );
FILL FILL_3_DFFPOSX1_4 ( );
FILL FILL_4_DFFPOSX1_4 ( );
FILL FILL_5_DFFPOSX1_4 ( );
FILL FILL_6_DFFPOSX1_4 ( );
FILL FILL_7_DFFPOSX1_4 ( );
FILL FILL_8_DFFPOSX1_4 ( );
FILL FILL_9_DFFPOSX1_4 ( );
FILL FILL_10_DFFPOSX1_4 ( );
FILL FILL_11_DFFPOSX1_4 ( );
FILL FILL_12_DFFPOSX1_4 ( );
FILL FILL_13_DFFPOSX1_4 ( );
FILL FILL_14_DFFPOSX1_4 ( );
FILL FILL_15_DFFPOSX1_4 ( );
FILL FILL_16_DFFPOSX1_4 ( );
FILL FILL_17_DFFPOSX1_4 ( );
FILL FILL_18_DFFPOSX1_4 ( );
FILL FILL_19_DFFPOSX1_4 ( );
FILL FILL_20_DFFPOSX1_4 ( );
FILL FILL_21_DFFPOSX1_4 ( );
FILL FILL_22_DFFPOSX1_4 ( );
FILL FILL_23_DFFPOSX1_4 ( );
FILL FILL_24_DFFPOSX1_4 ( );
FILL FILL_25_DFFPOSX1_4 ( );
FILL FILL_26_DFFPOSX1_4 ( );
FILL FILL_27_DFFPOSX1_4 ( );
FILL FILL_0_AND2X2_27 ( );
FILL FILL_1_AND2X2_27 ( );
FILL FILL_2_AND2X2_27 ( );
FILL FILL_3_AND2X2_27 ( );
FILL FILL_4_AND2X2_27 ( );
FILL FILL_5_AND2X2_27 ( );
FILL FILL_6_AND2X2_27 ( );
FILL FILL_7_AND2X2_27 ( );
FILL FILL_8_AND2X2_27 ( );
FILL FILL_0_NAND2X1_53 ( );
FILL FILL_1_NAND2X1_53 ( );
FILL FILL_2_NAND2X1_53 ( );
FILL FILL_3_NAND2X1_53 ( );
FILL FILL_4_NAND2X1_53 ( );
FILL FILL_5_NAND2X1_53 ( );
FILL FILL_6_NAND2X1_53 ( );
FILL FILL_0_NAND3X1_129 ( );
FILL FILL_1_NAND3X1_129 ( );
FILL FILL_2_NAND3X1_129 ( );
FILL FILL_3_NAND3X1_129 ( );
FILL FILL_4_NAND3X1_129 ( );
FILL FILL_5_NAND3X1_129 ( );
FILL FILL_6_NAND3X1_129 ( );
FILL FILL_7_NAND3X1_129 ( );
FILL FILL_8_NAND3X1_129 ( );
FILL FILL_0_AOI21X1_48 ( );
FILL FILL_1_AOI21X1_48 ( );
FILL FILL_2_AOI21X1_48 ( );
FILL FILL_3_AOI21X1_48 ( );
FILL FILL_4_AOI21X1_48 ( );
FILL FILL_5_AOI21X1_48 ( );
FILL FILL_6_AOI21X1_48 ( );
FILL FILL_7_AOI21X1_48 ( );
FILL FILL_8_AOI21X1_48 ( );
FILL FILL_0_INVX1_199 ( );
FILL FILL_1_INVX1_199 ( );
FILL FILL_2_INVX1_199 ( );
FILL FILL_3_INVX1_199 ( );
FILL FILL_4_INVX1_199 ( );
FILL FILL_0_DFFSR_62 ( );
FILL FILL_1_DFFSR_62 ( );
FILL FILL_2_DFFSR_62 ( );
FILL FILL_3_DFFSR_62 ( );
FILL FILL_4_DFFSR_62 ( );
FILL FILL_5_DFFSR_62 ( );
FILL FILL_6_DFFSR_62 ( );
FILL FILL_7_DFFSR_62 ( );
FILL FILL_8_DFFSR_62 ( );
FILL FILL_9_DFFSR_62 ( );
FILL FILL_10_DFFSR_62 ( );
FILL FILL_11_DFFSR_62 ( );
FILL FILL_12_DFFSR_62 ( );
FILL FILL_13_DFFSR_62 ( );
FILL FILL_14_DFFSR_62 ( );
FILL FILL_15_DFFSR_62 ( );
FILL FILL_16_DFFSR_62 ( );
FILL FILL_17_DFFSR_62 ( );
FILL FILL_18_DFFSR_62 ( );
FILL FILL_19_DFFSR_62 ( );
FILL FILL_20_DFFSR_62 ( );
FILL FILL_21_DFFSR_62 ( );
FILL FILL_22_DFFSR_62 ( );
FILL FILL_23_DFFSR_62 ( );
FILL FILL_24_DFFSR_62 ( );
FILL FILL_25_DFFSR_62 ( );
FILL FILL_26_DFFSR_62 ( );
FILL FILL_27_DFFSR_62 ( );
FILL FILL_28_DFFSR_62 ( );
FILL FILL_29_DFFSR_62 ( );
FILL FILL_30_DFFSR_62 ( );
FILL FILL_31_DFFSR_62 ( );
FILL FILL_32_DFFSR_62 ( );
FILL FILL_33_DFFSR_62 ( );
FILL FILL_34_DFFSR_62 ( );
FILL FILL_35_DFFSR_62 ( );
FILL FILL_36_DFFSR_62 ( );
FILL FILL_37_DFFSR_62 ( );
FILL FILL_38_DFFSR_62 ( );
FILL FILL_39_DFFSR_62 ( );
FILL FILL_40_DFFSR_62 ( );
FILL FILL_41_DFFSR_62 ( );
FILL FILL_42_DFFSR_62 ( );
FILL FILL_43_DFFSR_62 ( );
FILL FILL_44_DFFSR_62 ( );
FILL FILL_45_DFFSR_62 ( );
FILL FILL_46_DFFSR_62 ( );
FILL FILL_47_DFFSR_62 ( );
FILL FILL_48_DFFSR_62 ( );
FILL FILL_49_DFFSR_62 ( );
FILL FILL_50_DFFSR_62 ( );
FILL FILL_0_DFFSR_236 ( );
FILL FILL_1_DFFSR_236 ( );
FILL FILL_2_DFFSR_236 ( );
FILL FILL_3_DFFSR_236 ( );
FILL FILL_4_DFFSR_236 ( );
FILL FILL_5_DFFSR_236 ( );
FILL FILL_6_DFFSR_236 ( );
FILL FILL_7_DFFSR_236 ( );
FILL FILL_8_DFFSR_236 ( );
FILL FILL_9_DFFSR_236 ( );
FILL FILL_10_DFFSR_236 ( );
FILL FILL_11_DFFSR_236 ( );
FILL FILL_12_DFFSR_236 ( );
FILL FILL_13_DFFSR_236 ( );
FILL FILL_14_DFFSR_236 ( );
FILL FILL_15_DFFSR_236 ( );
FILL FILL_16_DFFSR_236 ( );
FILL FILL_17_DFFSR_236 ( );
FILL FILL_18_DFFSR_236 ( );
FILL FILL_19_DFFSR_236 ( );
FILL FILL_20_DFFSR_236 ( );
FILL FILL_21_DFFSR_236 ( );
FILL FILL_22_DFFSR_236 ( );
FILL FILL_23_DFFSR_236 ( );
FILL FILL_24_DFFSR_236 ( );
FILL FILL_25_DFFSR_236 ( );
FILL FILL_26_DFFSR_236 ( );
FILL FILL_27_DFFSR_236 ( );
FILL FILL_28_DFFSR_236 ( );
FILL FILL_29_DFFSR_236 ( );
FILL FILL_30_DFFSR_236 ( );
FILL FILL_31_DFFSR_236 ( );
FILL FILL_32_DFFSR_236 ( );
FILL FILL_33_DFFSR_236 ( );
FILL FILL_34_DFFSR_236 ( );
FILL FILL_35_DFFSR_236 ( );
FILL FILL_36_DFFSR_236 ( );
FILL FILL_37_DFFSR_236 ( );
FILL FILL_38_DFFSR_236 ( );
FILL FILL_39_DFFSR_236 ( );
FILL FILL_40_DFFSR_236 ( );
FILL FILL_41_DFFSR_236 ( );
FILL FILL_42_DFFSR_236 ( );
FILL FILL_43_DFFSR_236 ( );
FILL FILL_44_DFFSR_236 ( );
FILL FILL_45_DFFSR_236 ( );
FILL FILL_46_DFFSR_236 ( );
FILL FILL_47_DFFSR_236 ( );
FILL FILL_48_DFFSR_236 ( );
FILL FILL_49_DFFSR_236 ( );
FILL FILL_50_DFFSR_236 ( );
FILL FILL_0_NAND3X1_89 ( );
FILL FILL_1_NAND3X1_89 ( );
FILL FILL_2_NAND3X1_89 ( );
FILL FILL_3_NAND3X1_89 ( );
FILL FILL_4_NAND3X1_89 ( );
FILL FILL_5_NAND3X1_89 ( );
FILL FILL_6_NAND3X1_89 ( );
FILL FILL_7_NAND3X1_89 ( );
FILL FILL_8_NAND3X1_89 ( );
FILL FILL_0_NAND3X1_86 ( );
FILL FILL_1_NAND3X1_86 ( );
FILL FILL_2_NAND3X1_86 ( );
FILL FILL_3_NAND3X1_86 ( );
FILL FILL_4_NAND3X1_86 ( );
FILL FILL_5_NAND3X1_86 ( );
FILL FILL_6_NAND3X1_86 ( );
FILL FILL_7_NAND3X1_86 ( );
FILL FILL_8_NAND3X1_86 ( );
FILL FILL_0_INVX1_62 ( );
FILL FILL_1_INVX1_62 ( );
FILL FILL_2_INVX1_62 ( );
FILL FILL_3_INVX1_62 ( );
FILL FILL_0_DFFSR_169 ( );
FILL FILL_1_DFFSR_169 ( );
FILL FILL_2_DFFSR_169 ( );
FILL FILL_3_DFFSR_169 ( );
FILL FILL_4_DFFSR_169 ( );
FILL FILL_5_DFFSR_169 ( );
FILL FILL_6_DFFSR_169 ( );
FILL FILL_7_DFFSR_169 ( );
FILL FILL_8_DFFSR_169 ( );
FILL FILL_9_DFFSR_169 ( );
FILL FILL_10_DFFSR_169 ( );
FILL FILL_11_DFFSR_169 ( );
FILL FILL_12_DFFSR_169 ( );
FILL FILL_13_DFFSR_169 ( );
FILL FILL_14_DFFSR_169 ( );
FILL FILL_15_DFFSR_169 ( );
FILL FILL_16_DFFSR_169 ( );
FILL FILL_17_DFFSR_169 ( );
FILL FILL_18_DFFSR_169 ( );
FILL FILL_19_DFFSR_169 ( );
FILL FILL_20_DFFSR_169 ( );
FILL FILL_21_DFFSR_169 ( );
FILL FILL_22_DFFSR_169 ( );
FILL FILL_23_DFFSR_169 ( );
FILL FILL_24_DFFSR_169 ( );
FILL FILL_25_DFFSR_169 ( );
FILL FILL_26_DFFSR_169 ( );
FILL FILL_27_DFFSR_169 ( );
FILL FILL_28_DFFSR_169 ( );
FILL FILL_29_DFFSR_169 ( );
FILL FILL_30_DFFSR_169 ( );
FILL FILL_31_DFFSR_169 ( );
FILL FILL_32_DFFSR_169 ( );
FILL FILL_33_DFFSR_169 ( );
FILL FILL_34_DFFSR_169 ( );
FILL FILL_35_DFFSR_169 ( );
FILL FILL_36_DFFSR_169 ( );
FILL FILL_37_DFFSR_169 ( );
FILL FILL_38_DFFSR_169 ( );
FILL FILL_39_DFFSR_169 ( );
FILL FILL_40_DFFSR_169 ( );
FILL FILL_41_DFFSR_169 ( );
FILL FILL_42_DFFSR_169 ( );
FILL FILL_43_DFFSR_169 ( );
FILL FILL_44_DFFSR_169 ( );
FILL FILL_45_DFFSR_169 ( );
FILL FILL_46_DFFSR_169 ( );
FILL FILL_47_DFFSR_169 ( );
FILL FILL_48_DFFSR_169 ( );
FILL FILL_49_DFFSR_169 ( );
FILL FILL_50_DFFSR_169 ( );
FILL FILL_0_DFFSR_207 ( );
FILL FILL_1_DFFSR_207 ( );
FILL FILL_2_DFFSR_207 ( );
FILL FILL_3_DFFSR_207 ( );
FILL FILL_4_DFFSR_207 ( );
FILL FILL_5_DFFSR_207 ( );
FILL FILL_6_DFFSR_207 ( );
FILL FILL_7_DFFSR_207 ( );
FILL FILL_8_DFFSR_207 ( );
FILL FILL_9_DFFSR_207 ( );
FILL FILL_10_DFFSR_207 ( );
FILL FILL_11_DFFSR_207 ( );
FILL FILL_12_DFFSR_207 ( );
FILL FILL_13_DFFSR_207 ( );
FILL FILL_14_DFFSR_207 ( );
FILL FILL_15_DFFSR_207 ( );
FILL FILL_16_DFFSR_207 ( );
FILL FILL_17_DFFSR_207 ( );
FILL FILL_18_DFFSR_207 ( );
FILL FILL_19_DFFSR_207 ( );
FILL FILL_20_DFFSR_207 ( );
FILL FILL_21_DFFSR_207 ( );
FILL FILL_22_DFFSR_207 ( );
FILL FILL_23_DFFSR_207 ( );
FILL FILL_24_DFFSR_207 ( );
FILL FILL_25_DFFSR_207 ( );
FILL FILL_26_DFFSR_207 ( );
FILL FILL_27_DFFSR_207 ( );
FILL FILL_28_DFFSR_207 ( );
FILL FILL_29_DFFSR_207 ( );
FILL FILL_30_DFFSR_207 ( );
FILL FILL_31_DFFSR_207 ( );
FILL FILL_32_DFFSR_207 ( );
FILL FILL_33_DFFSR_207 ( );
FILL FILL_34_DFFSR_207 ( );
FILL FILL_35_DFFSR_207 ( );
FILL FILL_36_DFFSR_207 ( );
FILL FILL_37_DFFSR_207 ( );
FILL FILL_38_DFFSR_207 ( );
FILL FILL_39_DFFSR_207 ( );
FILL FILL_40_DFFSR_207 ( );
FILL FILL_41_DFFSR_207 ( );
FILL FILL_42_DFFSR_207 ( );
FILL FILL_43_DFFSR_207 ( );
FILL FILL_44_DFFSR_207 ( );
FILL FILL_45_DFFSR_207 ( );
FILL FILL_46_DFFSR_207 ( );
FILL FILL_47_DFFSR_207 ( );
FILL FILL_48_DFFSR_207 ( );
FILL FILL_49_DFFSR_207 ( );
FILL FILL_50_DFFSR_207 ( );
FILL FILL_0_NAND3X1_118 ( );
FILL FILL_1_NAND3X1_118 ( );
FILL FILL_2_NAND3X1_118 ( );
FILL FILL_3_NAND3X1_118 ( );
FILL FILL_4_NAND3X1_118 ( );
FILL FILL_5_NAND3X1_118 ( );
FILL FILL_6_NAND3X1_118 ( );
FILL FILL_7_NAND3X1_118 ( );
FILL FILL_8_NAND3X1_118 ( );
FILL FILL_0_NAND3X1_126 ( );
FILL FILL_1_NAND3X1_126 ( );
FILL FILL_2_NAND3X1_126 ( );
FILL FILL_3_NAND3X1_126 ( );
FILL FILL_4_NAND3X1_126 ( );
FILL FILL_5_NAND3X1_126 ( );
FILL FILL_6_NAND3X1_126 ( );
FILL FILL_7_NAND3X1_126 ( );
FILL FILL_8_NAND3X1_126 ( );
FILL FILL_9_NAND3X1_126 ( );
FILL FILL_0_NAND2X1_50 ( );
FILL FILL_1_NAND2X1_50 ( );
FILL FILL_2_NAND2X1_50 ( );
FILL FILL_3_NAND2X1_50 ( );
FILL FILL_4_NAND2X1_50 ( );
FILL FILL_5_NAND2X1_50 ( );
FILL FILL_6_NAND2X1_50 ( );
FILL FILL_0_DFFSR_200 ( );
FILL FILL_1_DFFSR_200 ( );
FILL FILL_2_DFFSR_200 ( );
FILL FILL_3_DFFSR_200 ( );
FILL FILL_4_DFFSR_200 ( );
FILL FILL_5_DFFSR_200 ( );
FILL FILL_6_DFFSR_200 ( );
FILL FILL_7_DFFSR_200 ( );
FILL FILL_8_DFFSR_200 ( );
FILL FILL_9_DFFSR_200 ( );
FILL FILL_10_DFFSR_200 ( );
FILL FILL_11_DFFSR_200 ( );
FILL FILL_12_DFFSR_200 ( );
FILL FILL_13_DFFSR_200 ( );
FILL FILL_14_DFFSR_200 ( );
FILL FILL_15_DFFSR_200 ( );
FILL FILL_16_DFFSR_200 ( );
FILL FILL_17_DFFSR_200 ( );
FILL FILL_18_DFFSR_200 ( );
FILL FILL_19_DFFSR_200 ( );
FILL FILL_20_DFFSR_200 ( );
FILL FILL_21_DFFSR_200 ( );
FILL FILL_22_DFFSR_200 ( );
FILL FILL_23_DFFSR_200 ( );
FILL FILL_24_DFFSR_200 ( );
FILL FILL_25_DFFSR_200 ( );
FILL FILL_26_DFFSR_200 ( );
FILL FILL_27_DFFSR_200 ( );
FILL FILL_28_DFFSR_200 ( );
FILL FILL_29_DFFSR_200 ( );
FILL FILL_30_DFFSR_200 ( );
FILL FILL_31_DFFSR_200 ( );
FILL FILL_32_DFFSR_200 ( );
FILL FILL_33_DFFSR_200 ( );
FILL FILL_34_DFFSR_200 ( );
FILL FILL_35_DFFSR_200 ( );
FILL FILL_36_DFFSR_200 ( );
FILL FILL_37_DFFSR_200 ( );
FILL FILL_38_DFFSR_200 ( );
FILL FILL_39_DFFSR_200 ( );
FILL FILL_40_DFFSR_200 ( );
FILL FILL_41_DFFSR_200 ( );
FILL FILL_42_DFFSR_200 ( );
FILL FILL_43_DFFSR_200 ( );
FILL FILL_44_DFFSR_200 ( );
FILL FILL_45_DFFSR_200 ( );
FILL FILL_46_DFFSR_200 ( );
FILL FILL_47_DFFSR_200 ( );
FILL FILL_48_DFFSR_200 ( );
FILL FILL_49_DFFSR_200 ( );
FILL FILL_50_DFFSR_200 ( );
FILL FILL_0_BUFX2_64 ( );
FILL FILL_1_BUFX2_64 ( );
FILL FILL_2_BUFX2_64 ( );
FILL FILL_3_BUFX2_64 ( );
FILL FILL_4_BUFX2_64 ( );
FILL FILL_5_BUFX2_64 ( );
FILL FILL_6_BUFX2_64 ( );
FILL FILL_0_AOI22X1_24 ( );
FILL FILL_1_AOI22X1_24 ( );
FILL FILL_2_AOI22X1_24 ( );
FILL FILL_3_AOI22X1_24 ( );
FILL FILL_4_AOI22X1_24 ( );
FILL FILL_5_AOI22X1_24 ( );
FILL FILL_6_AOI22X1_24 ( );
FILL FILL_7_AOI22X1_24 ( );
FILL FILL_8_AOI22X1_24 ( );
FILL FILL_9_AOI22X1_24 ( );
FILL FILL_10_AOI22X1_24 ( );
FILL FILL_11_AOI22X1_24 ( );
FILL FILL_0_NAND3X1_209 ( );
FILL FILL_1_NAND3X1_209 ( );
FILL FILL_2_NAND3X1_209 ( );
FILL FILL_3_NAND3X1_209 ( );
FILL FILL_4_NAND3X1_209 ( );
FILL FILL_5_NAND3X1_209 ( );
FILL FILL_6_NAND3X1_209 ( );
FILL FILL_7_NAND3X1_209 ( );
FILL FILL_8_NAND3X1_209 ( );
FILL FILL_0_NAND3X1_214 ( );
FILL FILL_1_NAND3X1_214 ( );
FILL FILL_2_NAND3X1_214 ( );
FILL FILL_3_NAND3X1_214 ( );
FILL FILL_4_NAND3X1_214 ( );
FILL FILL_5_NAND3X1_214 ( );
FILL FILL_6_NAND3X1_214 ( );
FILL FILL_7_NAND3X1_214 ( );
FILL FILL_8_NAND3X1_214 ( );
FILL FILL_9_NAND3X1_214 ( );
FILL FILL_0_NAND3X1_216 ( );
FILL FILL_1_NAND3X1_216 ( );
FILL FILL_2_NAND3X1_216 ( );
FILL FILL_3_NAND3X1_216 ( );
FILL FILL_4_NAND3X1_216 ( );
FILL FILL_5_NAND3X1_216 ( );
FILL FILL_6_NAND3X1_216 ( );
FILL FILL_7_NAND3X1_216 ( );
FILL FILL_8_NAND3X1_216 ( );
FILL FILL_0_DFFPOSX1_20 ( );
FILL FILL_1_DFFPOSX1_20 ( );
FILL FILL_2_DFFPOSX1_20 ( );
FILL FILL_3_DFFPOSX1_20 ( );
FILL FILL_4_DFFPOSX1_20 ( );
FILL FILL_5_DFFPOSX1_20 ( );
FILL FILL_6_DFFPOSX1_20 ( );
FILL FILL_7_DFFPOSX1_20 ( );
FILL FILL_8_DFFPOSX1_20 ( );
FILL FILL_9_DFFPOSX1_20 ( );
FILL FILL_10_DFFPOSX1_20 ( );
FILL FILL_11_DFFPOSX1_20 ( );
FILL FILL_12_DFFPOSX1_20 ( );
FILL FILL_13_DFFPOSX1_20 ( );
FILL FILL_14_DFFPOSX1_20 ( );
FILL FILL_15_DFFPOSX1_20 ( );
FILL FILL_16_DFFPOSX1_20 ( );
FILL FILL_17_DFFPOSX1_20 ( );
FILL FILL_18_DFFPOSX1_20 ( );
FILL FILL_19_DFFPOSX1_20 ( );
FILL FILL_20_DFFPOSX1_20 ( );
FILL FILL_21_DFFPOSX1_20 ( );
FILL FILL_22_DFFPOSX1_20 ( );
FILL FILL_23_DFFPOSX1_20 ( );
FILL FILL_24_DFFPOSX1_20 ( );
FILL FILL_25_DFFPOSX1_20 ( );
FILL FILL_26_DFFPOSX1_20 ( );
FILL FILL_27_DFFPOSX1_20 ( );
FILL FILL_0_NOR2X1_66 ( );
FILL FILL_1_NOR2X1_66 ( );
FILL FILL_2_NOR2X1_66 ( );
FILL FILL_3_NOR2X1_66 ( );
FILL FILL_4_NOR2X1_66 ( );
FILL FILL_5_NOR2X1_66 ( );
FILL FILL_6_NOR2X1_66 ( );
FILL FILL_0_NAND3X1_141 ( );
FILL FILL_1_NAND3X1_141 ( );
FILL FILL_2_NAND3X1_141 ( );
FILL FILL_3_NAND3X1_141 ( );
FILL FILL_4_NAND3X1_141 ( );
FILL FILL_5_NAND3X1_141 ( );
FILL FILL_6_NAND3X1_141 ( );
FILL FILL_7_NAND3X1_141 ( );
FILL FILL_8_NAND3X1_141 ( );
FILL FILL_0_NAND2X1_64 ( );
FILL FILL_1_NAND2X1_64 ( );
FILL FILL_2_NAND2X1_64 ( );
FILL FILL_3_NAND2X1_64 ( );
FILL FILL_4_NAND2X1_64 ( );
FILL FILL_5_NAND2X1_64 ( );
FILL FILL_6_NAND2X1_64 ( );
FILL FILL_0_NAND3X1_195 ( );
FILL FILL_1_NAND3X1_195 ( );
FILL FILL_2_NAND3X1_195 ( );
FILL FILL_3_NAND3X1_195 ( );
FILL FILL_4_NAND3X1_195 ( );
FILL FILL_5_NAND3X1_195 ( );
FILL FILL_6_NAND3X1_195 ( );
FILL FILL_7_NAND3X1_195 ( );
FILL FILL_8_NAND3X1_195 ( );
FILL FILL_0_OAI21X1_74 ( );
FILL FILL_1_OAI21X1_74 ( );
FILL FILL_2_OAI21X1_74 ( );
FILL FILL_3_OAI21X1_74 ( );
FILL FILL_4_OAI21X1_74 ( );
FILL FILL_5_OAI21X1_74 ( );
FILL FILL_6_OAI21X1_74 ( );
FILL FILL_7_OAI21X1_74 ( );
FILL FILL_8_OAI21X1_74 ( );
FILL FILL_0_NAND3X1_196 ( );
FILL FILL_1_NAND3X1_196 ( );
FILL FILL_2_NAND3X1_196 ( );
FILL FILL_3_NAND3X1_196 ( );
FILL FILL_4_NAND3X1_196 ( );
FILL FILL_5_NAND3X1_196 ( );
FILL FILL_6_NAND3X1_196 ( );
FILL FILL_7_NAND3X1_196 ( );
FILL FILL_8_NAND3X1_196 ( );
FILL FILL_0_DFFPOSX1_18 ( );
FILL FILL_1_DFFPOSX1_18 ( );
FILL FILL_2_DFFPOSX1_18 ( );
FILL FILL_3_DFFPOSX1_18 ( );
FILL FILL_4_DFFPOSX1_18 ( );
FILL FILL_5_DFFPOSX1_18 ( );
FILL FILL_6_DFFPOSX1_18 ( );
FILL FILL_7_DFFPOSX1_18 ( );
FILL FILL_8_DFFPOSX1_18 ( );
FILL FILL_9_DFFPOSX1_18 ( );
FILL FILL_10_DFFPOSX1_18 ( );
FILL FILL_11_DFFPOSX1_18 ( );
FILL FILL_12_DFFPOSX1_18 ( );
FILL FILL_13_DFFPOSX1_18 ( );
FILL FILL_14_DFFPOSX1_18 ( );
FILL FILL_15_DFFPOSX1_18 ( );
FILL FILL_16_DFFPOSX1_18 ( );
FILL FILL_17_DFFPOSX1_18 ( );
FILL FILL_18_DFFPOSX1_18 ( );
FILL FILL_19_DFFPOSX1_18 ( );
FILL FILL_20_DFFPOSX1_18 ( );
FILL FILL_21_DFFPOSX1_18 ( );
FILL FILL_22_DFFPOSX1_18 ( );
FILL FILL_23_DFFPOSX1_18 ( );
FILL FILL_24_DFFPOSX1_18 ( );
FILL FILL_25_DFFPOSX1_18 ( );
FILL FILL_26_DFFPOSX1_18 ( );
FILL FILL_27_DFFPOSX1_18 ( );
FILL FILL_0_OAI21X1_17 ( );
FILL FILL_1_OAI21X1_17 ( );
FILL FILL_2_OAI21X1_17 ( );
FILL FILL_3_OAI21X1_17 ( );
FILL FILL_4_OAI21X1_17 ( );
FILL FILL_5_OAI21X1_17 ( );
FILL FILL_6_OAI21X1_17 ( );
FILL FILL_7_OAI21X1_17 ( );
FILL FILL_8_OAI21X1_17 ( );
FILL FILL_0_NAND2X1_144 ( );
FILL FILL_1_NAND2X1_144 ( );
FILL FILL_2_NAND2X1_144 ( );
FILL FILL_3_NAND2X1_144 ( );
FILL FILL_4_NAND2X1_144 ( );
FILL FILL_5_NAND2X1_144 ( );
FILL FILL_6_NAND2X1_144 ( );
FILL FILL_0_NAND2X1_141 ( );
FILL FILL_1_NAND2X1_141 ( );
FILL FILL_2_NAND2X1_141 ( );
FILL FILL_3_NAND2X1_141 ( );
FILL FILL_4_NAND2X1_141 ( );
FILL FILL_5_NAND2X1_141 ( );
FILL FILL_6_NAND2X1_141 ( );
FILL FILL_0_CLKBUF1_15 ( );
FILL FILL_1_CLKBUF1_15 ( );
FILL FILL_2_CLKBUF1_15 ( );
FILL FILL_3_CLKBUF1_15 ( );
FILL FILL_4_CLKBUF1_15 ( );
FILL FILL_5_CLKBUF1_15 ( );
FILL FILL_6_CLKBUF1_15 ( );
FILL FILL_7_CLKBUF1_15 ( );
FILL FILL_8_CLKBUF1_15 ( );
FILL FILL_9_CLKBUF1_15 ( );
FILL FILL_10_CLKBUF1_15 ( );
FILL FILL_11_CLKBUF1_15 ( );
FILL FILL_12_CLKBUF1_15 ( );
FILL FILL_13_CLKBUF1_15 ( );
FILL FILL_14_CLKBUF1_15 ( );
FILL FILL_15_CLKBUF1_15 ( );
FILL FILL_16_CLKBUF1_15 ( );
FILL FILL_17_CLKBUF1_15 ( );
FILL FILL_18_CLKBUF1_15 ( );
FILL FILL_19_CLKBUF1_15 ( );
FILL FILL_20_CLKBUF1_15 ( );
FILL FILL_0_INVX1_97 ( );
FILL FILL_1_INVX1_97 ( );
FILL FILL_2_INVX1_97 ( );
FILL FILL_3_INVX1_97 ( );
FILL FILL_4_INVX1_97 ( );
FILL FILL_0_DFFSR_172 ( );
FILL FILL_1_DFFSR_172 ( );
FILL FILL_2_DFFSR_172 ( );
FILL FILL_3_DFFSR_172 ( );
FILL FILL_4_DFFSR_172 ( );
FILL FILL_5_DFFSR_172 ( );
FILL FILL_6_DFFSR_172 ( );
FILL FILL_7_DFFSR_172 ( );
FILL FILL_8_DFFSR_172 ( );
FILL FILL_9_DFFSR_172 ( );
FILL FILL_10_DFFSR_172 ( );
FILL FILL_11_DFFSR_172 ( );
FILL FILL_12_DFFSR_172 ( );
FILL FILL_13_DFFSR_172 ( );
FILL FILL_14_DFFSR_172 ( );
FILL FILL_15_DFFSR_172 ( );
FILL FILL_16_DFFSR_172 ( );
FILL FILL_17_DFFSR_172 ( );
FILL FILL_18_DFFSR_172 ( );
FILL FILL_19_DFFSR_172 ( );
FILL FILL_20_DFFSR_172 ( );
FILL FILL_21_DFFSR_172 ( );
FILL FILL_22_DFFSR_172 ( );
FILL FILL_23_DFFSR_172 ( );
FILL FILL_24_DFFSR_172 ( );
FILL FILL_25_DFFSR_172 ( );
FILL FILL_26_DFFSR_172 ( );
FILL FILL_27_DFFSR_172 ( );
FILL FILL_28_DFFSR_172 ( );
FILL FILL_29_DFFSR_172 ( );
FILL FILL_30_DFFSR_172 ( );
FILL FILL_31_DFFSR_172 ( );
FILL FILL_32_DFFSR_172 ( );
FILL FILL_33_DFFSR_172 ( );
FILL FILL_34_DFFSR_172 ( );
FILL FILL_35_DFFSR_172 ( );
FILL FILL_36_DFFSR_172 ( );
FILL FILL_37_DFFSR_172 ( );
FILL FILL_38_DFFSR_172 ( );
FILL FILL_39_DFFSR_172 ( );
FILL FILL_40_DFFSR_172 ( );
FILL FILL_41_DFFSR_172 ( );
FILL FILL_42_DFFSR_172 ( );
FILL FILL_43_DFFSR_172 ( );
FILL FILL_44_DFFSR_172 ( );
FILL FILL_45_DFFSR_172 ( );
FILL FILL_46_DFFSR_172 ( );
FILL FILL_47_DFFSR_172 ( );
FILL FILL_48_DFFSR_172 ( );
FILL FILL_49_DFFSR_172 ( );
FILL FILL_50_DFFSR_172 ( );
FILL FILL_0_INVX1_99 ( );
FILL FILL_1_INVX1_99 ( );
FILL FILL_2_INVX1_99 ( );
FILL FILL_3_INVX1_99 ( );
FILL FILL_4_INVX1_99 ( );
FILL FILL_0_NAND2X1_116 ( );
FILL FILL_1_NAND2X1_116 ( );
FILL FILL_2_NAND2X1_116 ( );
FILL FILL_3_NAND2X1_116 ( );
FILL FILL_4_NAND2X1_116 ( );
FILL FILL_5_NAND2X1_116 ( );
FILL FILL_6_NAND2X1_116 ( );
FILL FILL_0_INVX1_78 ( );
FILL FILL_1_INVX1_78 ( );
FILL FILL_2_INVX1_78 ( );
FILL FILL_3_INVX1_78 ( );
FILL FILL_4_INVX1_78 ( );
FILL FILL_0_INVX1_98 ( );
FILL FILL_1_INVX1_98 ( );
FILL FILL_2_INVX1_98 ( );
FILL FILL_3_INVX1_98 ( );
FILL FILL_0_OAI22X1_40 ( );
FILL FILL_1_OAI22X1_40 ( );
FILL FILL_2_OAI22X1_40 ( );
FILL FILL_3_OAI22X1_40 ( );
FILL FILL_4_OAI22X1_40 ( );
FILL FILL_5_OAI22X1_40 ( );
FILL FILL_6_OAI22X1_40 ( );
FILL FILL_7_OAI22X1_40 ( );
FILL FILL_8_OAI22X1_40 ( );
FILL FILL_9_OAI22X1_40 ( );
FILL FILL_10_OAI22X1_40 ( );
FILL FILL_11_OAI22X1_40 ( );
FILL FILL_0_NAND3X1_87 ( );
FILL FILL_1_NAND3X1_87 ( );
FILL FILL_2_NAND3X1_87 ( );
FILL FILL_3_NAND3X1_87 ( );
FILL FILL_4_NAND3X1_87 ( );
FILL FILL_5_NAND3X1_87 ( );
FILL FILL_6_NAND3X1_87 ( );
FILL FILL_7_NAND3X1_87 ( );
FILL FILL_8_NAND3X1_87 ( );
FILL FILL_0_NAND3X1_85 ( );
FILL FILL_1_NAND3X1_85 ( );
FILL FILL_2_NAND3X1_85 ( );
FILL FILL_3_NAND3X1_85 ( );
FILL FILL_4_NAND3X1_85 ( );
FILL FILL_5_NAND3X1_85 ( );
FILL FILL_6_NAND3X1_85 ( );
FILL FILL_7_NAND3X1_85 ( );
FILL FILL_8_NAND3X1_85 ( );
FILL FILL_0_DFFSR_195 ( );
FILL FILL_1_DFFSR_195 ( );
FILL FILL_2_DFFSR_195 ( );
FILL FILL_3_DFFSR_195 ( );
FILL FILL_4_DFFSR_195 ( );
FILL FILL_5_DFFSR_195 ( );
FILL FILL_6_DFFSR_195 ( );
FILL FILL_7_DFFSR_195 ( );
FILL FILL_8_DFFSR_195 ( );
FILL FILL_9_DFFSR_195 ( );
FILL FILL_10_DFFSR_195 ( );
FILL FILL_11_DFFSR_195 ( );
FILL FILL_12_DFFSR_195 ( );
FILL FILL_13_DFFSR_195 ( );
FILL FILL_14_DFFSR_195 ( );
FILL FILL_15_DFFSR_195 ( );
FILL FILL_16_DFFSR_195 ( );
FILL FILL_17_DFFSR_195 ( );
FILL FILL_18_DFFSR_195 ( );
FILL FILL_19_DFFSR_195 ( );
FILL FILL_20_DFFSR_195 ( );
FILL FILL_21_DFFSR_195 ( );
FILL FILL_22_DFFSR_195 ( );
FILL FILL_23_DFFSR_195 ( );
FILL FILL_24_DFFSR_195 ( );
FILL FILL_25_DFFSR_195 ( );
FILL FILL_26_DFFSR_195 ( );
FILL FILL_27_DFFSR_195 ( );
FILL FILL_28_DFFSR_195 ( );
FILL FILL_29_DFFSR_195 ( );
FILL FILL_30_DFFSR_195 ( );
FILL FILL_31_DFFSR_195 ( );
FILL FILL_32_DFFSR_195 ( );
FILL FILL_33_DFFSR_195 ( );
FILL FILL_34_DFFSR_195 ( );
FILL FILL_35_DFFSR_195 ( );
FILL FILL_36_DFFSR_195 ( );
FILL FILL_37_DFFSR_195 ( );
FILL FILL_38_DFFSR_195 ( );
FILL FILL_39_DFFSR_195 ( );
FILL FILL_40_DFFSR_195 ( );
FILL FILL_41_DFFSR_195 ( );
FILL FILL_42_DFFSR_195 ( );
FILL FILL_43_DFFSR_195 ( );
FILL FILL_44_DFFSR_195 ( );
FILL FILL_45_DFFSR_195 ( );
FILL FILL_46_DFFSR_195 ( );
FILL FILL_47_DFFSR_195 ( );
FILL FILL_48_DFFSR_195 ( );
FILL FILL_49_DFFSR_195 ( );
FILL FILL_50_DFFSR_195 ( );
FILL FILL_0_BUFX2_28 ( );
FILL FILL_1_BUFX2_28 ( );
FILL FILL_2_BUFX2_28 ( );
FILL FILL_3_BUFX2_28 ( );
FILL FILL_4_BUFX2_28 ( );
FILL FILL_5_BUFX2_28 ( );
FILL FILL_6_BUFX2_28 ( );
FILL FILL_0_DFFSR_231 ( );
FILL FILL_1_DFFSR_231 ( );
FILL FILL_2_DFFSR_231 ( );
FILL FILL_3_DFFSR_231 ( );
FILL FILL_4_DFFSR_231 ( );
FILL FILL_5_DFFSR_231 ( );
FILL FILL_6_DFFSR_231 ( );
FILL FILL_7_DFFSR_231 ( );
FILL FILL_8_DFFSR_231 ( );
FILL FILL_9_DFFSR_231 ( );
FILL FILL_10_DFFSR_231 ( );
FILL FILL_11_DFFSR_231 ( );
FILL FILL_12_DFFSR_231 ( );
FILL FILL_13_DFFSR_231 ( );
FILL FILL_14_DFFSR_231 ( );
FILL FILL_15_DFFSR_231 ( );
FILL FILL_16_DFFSR_231 ( );
FILL FILL_17_DFFSR_231 ( );
FILL FILL_18_DFFSR_231 ( );
FILL FILL_19_DFFSR_231 ( );
FILL FILL_20_DFFSR_231 ( );
FILL FILL_21_DFFSR_231 ( );
FILL FILL_22_DFFSR_231 ( );
FILL FILL_23_DFFSR_231 ( );
FILL FILL_24_DFFSR_231 ( );
FILL FILL_25_DFFSR_231 ( );
FILL FILL_26_DFFSR_231 ( );
FILL FILL_27_DFFSR_231 ( );
FILL FILL_28_DFFSR_231 ( );
FILL FILL_29_DFFSR_231 ( );
FILL FILL_30_DFFSR_231 ( );
FILL FILL_31_DFFSR_231 ( );
FILL FILL_32_DFFSR_231 ( );
FILL FILL_33_DFFSR_231 ( );
FILL FILL_34_DFFSR_231 ( );
FILL FILL_35_DFFSR_231 ( );
FILL FILL_36_DFFSR_231 ( );
FILL FILL_37_DFFSR_231 ( );
FILL FILL_38_DFFSR_231 ( );
FILL FILL_39_DFFSR_231 ( );
FILL FILL_40_DFFSR_231 ( );
FILL FILL_41_DFFSR_231 ( );
FILL FILL_42_DFFSR_231 ( );
FILL FILL_43_DFFSR_231 ( );
FILL FILL_44_DFFSR_231 ( );
FILL FILL_45_DFFSR_231 ( );
FILL FILL_46_DFFSR_231 ( );
FILL FILL_47_DFFSR_231 ( );
FILL FILL_48_DFFSR_231 ( );
FILL FILL_49_DFFSR_231 ( );
FILL FILL_50_DFFSR_231 ( );
FILL FILL_0_NAND3X1_127 ( );
FILL FILL_1_NAND3X1_127 ( );
FILL FILL_2_NAND3X1_127 ( );
FILL FILL_3_NAND3X1_127 ( );
FILL FILL_4_NAND3X1_127 ( );
FILL FILL_5_NAND3X1_127 ( );
FILL FILL_6_NAND3X1_127 ( );
FILL FILL_7_NAND3X1_127 ( );
FILL FILL_8_NAND3X1_127 ( );
FILL FILL_9_NAND3X1_127 ( );
FILL FILL_0_INVX1_64 ( );
FILL FILL_1_INVX1_64 ( );
FILL FILL_2_INVX1_64 ( );
FILL FILL_3_INVX1_64 ( );
FILL FILL_4_INVX1_64 ( );
FILL FILL_0_BUFX2_62 ( );
FILL FILL_1_BUFX2_62 ( );
FILL FILL_2_BUFX2_62 ( );
FILL FILL_3_BUFX2_62 ( );
FILL FILL_4_BUFX2_62 ( );
FILL FILL_5_BUFX2_62 ( );
FILL FILL_6_BUFX2_62 ( );
FILL FILL_0_DFFSR_144 ( );
FILL FILL_1_DFFSR_144 ( );
FILL FILL_2_DFFSR_144 ( );
FILL FILL_3_DFFSR_144 ( );
FILL FILL_4_DFFSR_144 ( );
FILL FILL_5_DFFSR_144 ( );
FILL FILL_6_DFFSR_144 ( );
FILL FILL_7_DFFSR_144 ( );
FILL FILL_8_DFFSR_144 ( );
FILL FILL_9_DFFSR_144 ( );
FILL FILL_10_DFFSR_144 ( );
FILL FILL_11_DFFSR_144 ( );
FILL FILL_12_DFFSR_144 ( );
FILL FILL_13_DFFSR_144 ( );
FILL FILL_14_DFFSR_144 ( );
FILL FILL_15_DFFSR_144 ( );
FILL FILL_16_DFFSR_144 ( );
FILL FILL_17_DFFSR_144 ( );
FILL FILL_18_DFFSR_144 ( );
FILL FILL_19_DFFSR_144 ( );
FILL FILL_20_DFFSR_144 ( );
FILL FILL_21_DFFSR_144 ( );
FILL FILL_22_DFFSR_144 ( );
FILL FILL_23_DFFSR_144 ( );
FILL FILL_24_DFFSR_144 ( );
FILL FILL_25_DFFSR_144 ( );
FILL FILL_26_DFFSR_144 ( );
FILL FILL_27_DFFSR_144 ( );
FILL FILL_28_DFFSR_144 ( );
FILL FILL_29_DFFSR_144 ( );
FILL FILL_30_DFFSR_144 ( );
FILL FILL_31_DFFSR_144 ( );
FILL FILL_32_DFFSR_144 ( );
FILL FILL_33_DFFSR_144 ( );
FILL FILL_34_DFFSR_144 ( );
FILL FILL_35_DFFSR_144 ( );
FILL FILL_36_DFFSR_144 ( );
FILL FILL_37_DFFSR_144 ( );
FILL FILL_38_DFFSR_144 ( );
FILL FILL_39_DFFSR_144 ( );
FILL FILL_40_DFFSR_144 ( );
FILL FILL_41_DFFSR_144 ( );
FILL FILL_42_DFFSR_144 ( );
FILL FILL_43_DFFSR_144 ( );
FILL FILL_44_DFFSR_144 ( );
FILL FILL_45_DFFSR_144 ( );
FILL FILL_46_DFFSR_144 ( );
FILL FILL_47_DFFSR_144 ( );
FILL FILL_48_DFFSR_144 ( );
FILL FILL_49_DFFSR_144 ( );
FILL FILL_50_DFFSR_144 ( );
FILL FILL_0_NAND2X1_89 ( );
FILL FILL_1_NAND2X1_89 ( );
FILL FILL_2_NAND2X1_89 ( );
FILL FILL_3_NAND2X1_89 ( );
FILL FILL_4_NAND2X1_89 ( );
FILL FILL_5_NAND2X1_89 ( );
FILL FILL_6_NAND2X1_89 ( );
FILL FILL_0_OAI21X1_73 ( );
FILL FILL_1_OAI21X1_73 ( );
FILL FILL_2_OAI21X1_73 ( );
FILL FILL_3_OAI21X1_73 ( );
FILL FILL_4_OAI21X1_73 ( );
FILL FILL_5_OAI21X1_73 ( );
FILL FILL_6_OAI21X1_73 ( );
FILL FILL_7_OAI21X1_73 ( );
FILL FILL_8_OAI21X1_73 ( );
FILL FILL_0_NAND3X1_208 ( );
FILL FILL_1_NAND3X1_208 ( );
FILL FILL_2_NAND3X1_208 ( );
FILL FILL_3_NAND3X1_208 ( );
FILL FILL_4_NAND3X1_208 ( );
FILL FILL_5_NAND3X1_208 ( );
FILL FILL_6_NAND3X1_208 ( );
FILL FILL_7_NAND3X1_208 ( );
FILL FILL_8_NAND3X1_208 ( );
FILL FILL_9_NAND3X1_208 ( );
FILL FILL_0_NAND3X1_218 ( );
FILL FILL_1_NAND3X1_218 ( );
FILL FILL_2_NAND3X1_218 ( );
FILL FILL_3_NAND3X1_218 ( );
FILL FILL_4_NAND3X1_218 ( );
FILL FILL_5_NAND3X1_218 ( );
FILL FILL_6_NAND3X1_218 ( );
FILL FILL_7_NAND3X1_218 ( );
FILL FILL_8_NAND3X1_218 ( );
FILL FILL_0_NAND3X1_217 ( );
FILL FILL_1_NAND3X1_217 ( );
FILL FILL_2_NAND3X1_217 ( );
FILL FILL_3_NAND3X1_217 ( );
FILL FILL_4_NAND3X1_217 ( );
FILL FILL_5_NAND3X1_217 ( );
FILL FILL_6_NAND3X1_217 ( );
FILL FILL_7_NAND3X1_217 ( );
FILL FILL_8_NAND3X1_217 ( );
FILL FILL_9_NAND3X1_217 ( );
FILL FILL_0_NAND3X1_222 ( );
FILL FILL_1_NAND3X1_222 ( );
FILL FILL_2_NAND3X1_222 ( );
FILL FILL_3_NAND3X1_222 ( );
FILL FILL_4_NAND3X1_222 ( );
FILL FILL_5_NAND3X1_222 ( );
FILL FILL_6_NAND3X1_222 ( );
FILL FILL_7_NAND3X1_222 ( );
FILL FILL_8_NAND3X1_222 ( );
FILL FILL_0_NAND3X1_223 ( );
FILL FILL_1_NAND3X1_223 ( );
FILL FILL_2_NAND3X1_223 ( );
FILL FILL_3_NAND3X1_223 ( );
FILL FILL_4_NAND3X1_223 ( );
FILL FILL_5_NAND3X1_223 ( );
FILL FILL_6_NAND3X1_223 ( );
FILL FILL_7_NAND3X1_223 ( );
FILL FILL_8_NAND3X1_223 ( );
FILL FILL_9_NAND3X1_223 ( );
FILL FILL_0_NAND3X1_220 ( );
FILL FILL_1_NAND3X1_220 ( );
FILL FILL_2_NAND3X1_220 ( );
FILL FILL_3_NAND3X1_220 ( );
FILL FILL_4_NAND3X1_220 ( );
FILL FILL_5_NAND3X1_220 ( );
FILL FILL_6_NAND3X1_220 ( );
FILL FILL_7_NAND3X1_220 ( );
FILL FILL_8_NAND3X1_220 ( );
FILL FILL_9_NAND3X1_220 ( );
FILL FILL_0_NAND3X1_221 ( );
FILL FILL_1_NAND3X1_221 ( );
FILL FILL_2_NAND3X1_221 ( );
FILL FILL_3_NAND3X1_221 ( );
FILL FILL_4_NAND3X1_221 ( );
FILL FILL_5_NAND3X1_221 ( );
FILL FILL_6_NAND3X1_221 ( );
FILL FILL_7_NAND3X1_221 ( );
FILL FILL_8_NAND3X1_221 ( );
FILL FILL_0_NAND2X1_90 ( );
FILL FILL_1_NAND2X1_90 ( );
FILL FILL_2_NAND2X1_90 ( );
FILL FILL_3_NAND2X1_90 ( );
FILL FILL_4_NAND2X1_90 ( );
FILL FILL_5_NAND2X1_90 ( );
FILL FILL_6_NAND2X1_90 ( );
FILL FILL_0_AOI21X1_24 ( );
FILL FILL_1_AOI21X1_24 ( );
FILL FILL_2_AOI21X1_24 ( );
FILL FILL_3_AOI21X1_24 ( );
FILL FILL_4_AOI21X1_24 ( );
FILL FILL_5_AOI21X1_24 ( );
FILL FILL_6_AOI21X1_24 ( );
FILL FILL_7_AOI21X1_24 ( );
FILL FILL_8_AOI21X1_24 ( );
FILL FILL_9_AOI21X1_24 ( );
FILL FILL_0_OAI21X1_56 ( );
FILL FILL_1_OAI21X1_56 ( );
FILL FILL_2_OAI21X1_56 ( );
FILL FILL_3_OAI21X1_56 ( );
FILL FILL_4_OAI21X1_56 ( );
FILL FILL_5_OAI21X1_56 ( );
FILL FILL_6_OAI21X1_56 ( );
FILL FILL_7_OAI21X1_56 ( );
FILL FILL_8_OAI21X1_56 ( );
FILL FILL_0_NAND3X1_197 ( );
FILL FILL_1_NAND3X1_197 ( );
FILL FILL_2_NAND3X1_197 ( );
FILL FILL_3_NAND3X1_197 ( );
FILL FILL_4_NAND3X1_197 ( );
FILL FILL_5_NAND3X1_197 ( );
FILL FILL_6_NAND3X1_197 ( );
FILL FILL_7_NAND3X1_197 ( );
FILL FILL_8_NAND3X1_197 ( );
FILL FILL_0_NAND2X1_129 ( );
FILL FILL_1_NAND2X1_129 ( );
FILL FILL_2_NAND2X1_129 ( );
FILL FILL_3_NAND2X1_129 ( );
FILL FILL_4_NAND2X1_129 ( );
FILL FILL_5_NAND2X1_129 ( );
FILL FILL_6_NAND2X1_129 ( );
FILL FILL_0_OAI21X1_98 ( );
FILL FILL_1_OAI21X1_98 ( );
FILL FILL_2_OAI21X1_98 ( );
FILL FILL_3_OAI21X1_98 ( );
FILL FILL_4_OAI21X1_98 ( );
FILL FILL_5_OAI21X1_98 ( );
FILL FILL_6_OAI21X1_98 ( );
FILL FILL_7_OAI21X1_98 ( );
FILL FILL_8_OAI21X1_98 ( );
FILL FILL_9_OAI21X1_98 ( );
FILL FILL_0_INVX1_195 ( );
FILL FILL_1_INVX1_195 ( );
FILL FILL_2_INVX1_195 ( );
FILL FILL_3_INVX1_195 ( );
FILL FILL_0_NOR2X1_79 ( );
FILL FILL_1_NOR2X1_79 ( );
FILL FILL_2_NOR2X1_79 ( );
FILL FILL_3_NOR2X1_79 ( );
FILL FILL_4_NOR2X1_79 ( );
FILL FILL_5_NOR2X1_79 ( );
FILL FILL_6_NOR2X1_79 ( );
FILL FILL_0_INVX1_119 ( );
FILL FILL_1_INVX1_119 ( );
FILL FILL_2_INVX1_119 ( );
FILL FILL_3_INVX1_119 ( );
FILL FILL_4_INVX1_119 ( );
FILL FILL_0_DFFSR_46 ( );
FILL FILL_1_DFFSR_46 ( );
FILL FILL_2_DFFSR_46 ( );
FILL FILL_3_DFFSR_46 ( );
FILL FILL_4_DFFSR_46 ( );
FILL FILL_5_DFFSR_46 ( );
FILL FILL_6_DFFSR_46 ( );
FILL FILL_7_DFFSR_46 ( );
FILL FILL_8_DFFSR_46 ( );
FILL FILL_9_DFFSR_46 ( );
FILL FILL_10_DFFSR_46 ( );
FILL FILL_11_DFFSR_46 ( );
FILL FILL_12_DFFSR_46 ( );
FILL FILL_13_DFFSR_46 ( );
FILL FILL_14_DFFSR_46 ( );
FILL FILL_15_DFFSR_46 ( );
FILL FILL_16_DFFSR_46 ( );
FILL FILL_17_DFFSR_46 ( );
FILL FILL_18_DFFSR_46 ( );
FILL FILL_19_DFFSR_46 ( );
FILL FILL_20_DFFSR_46 ( );
FILL FILL_21_DFFSR_46 ( );
FILL FILL_22_DFFSR_46 ( );
FILL FILL_23_DFFSR_46 ( );
FILL FILL_24_DFFSR_46 ( );
FILL FILL_25_DFFSR_46 ( );
FILL FILL_26_DFFSR_46 ( );
FILL FILL_27_DFFSR_46 ( );
FILL FILL_28_DFFSR_46 ( );
FILL FILL_29_DFFSR_46 ( );
FILL FILL_30_DFFSR_46 ( );
FILL FILL_31_DFFSR_46 ( );
FILL FILL_32_DFFSR_46 ( );
FILL FILL_33_DFFSR_46 ( );
FILL FILL_34_DFFSR_46 ( );
FILL FILL_35_DFFSR_46 ( );
FILL FILL_36_DFFSR_46 ( );
FILL FILL_37_DFFSR_46 ( );
FILL FILL_38_DFFSR_46 ( );
FILL FILL_39_DFFSR_46 ( );
FILL FILL_40_DFFSR_46 ( );
FILL FILL_41_DFFSR_46 ( );
FILL FILL_42_DFFSR_46 ( );
FILL FILL_43_DFFSR_46 ( );
FILL FILL_44_DFFSR_46 ( );
FILL FILL_45_DFFSR_46 ( );
FILL FILL_46_DFFSR_46 ( );
FILL FILL_47_DFFSR_46 ( );
FILL FILL_48_DFFSR_46 ( );
FILL FILL_49_DFFSR_46 ( );
FILL FILL_50_DFFSR_46 ( );
FILL FILL_0_INVX1_86 ( );
FILL FILL_1_INVX1_86 ( );
FILL FILL_2_INVX1_86 ( );
FILL FILL_3_INVX1_86 ( );
FILL FILL_4_INVX1_86 ( );
FILL FILL_0_INVX1_85 ( );
FILL FILL_1_INVX1_85 ( );
FILL FILL_2_INVX1_85 ( );
FILL FILL_3_INVX1_85 ( );
FILL FILL_0_DFFSR_188 ( );
FILL FILL_1_DFFSR_188 ( );
FILL FILL_2_DFFSR_188 ( );
FILL FILL_3_DFFSR_188 ( );
FILL FILL_4_DFFSR_188 ( );
FILL FILL_5_DFFSR_188 ( );
FILL FILL_6_DFFSR_188 ( );
FILL FILL_7_DFFSR_188 ( );
FILL FILL_8_DFFSR_188 ( );
FILL FILL_9_DFFSR_188 ( );
FILL FILL_10_DFFSR_188 ( );
FILL FILL_11_DFFSR_188 ( );
FILL FILL_12_DFFSR_188 ( );
FILL FILL_13_DFFSR_188 ( );
FILL FILL_14_DFFSR_188 ( );
FILL FILL_15_DFFSR_188 ( );
FILL FILL_16_DFFSR_188 ( );
FILL FILL_17_DFFSR_188 ( );
FILL FILL_18_DFFSR_188 ( );
FILL FILL_19_DFFSR_188 ( );
FILL FILL_20_DFFSR_188 ( );
FILL FILL_21_DFFSR_188 ( );
FILL FILL_22_DFFSR_188 ( );
FILL FILL_23_DFFSR_188 ( );
FILL FILL_24_DFFSR_188 ( );
FILL FILL_25_DFFSR_188 ( );
FILL FILL_26_DFFSR_188 ( );
FILL FILL_27_DFFSR_188 ( );
FILL FILL_28_DFFSR_188 ( );
FILL FILL_29_DFFSR_188 ( );
FILL FILL_30_DFFSR_188 ( );
FILL FILL_31_DFFSR_188 ( );
FILL FILL_32_DFFSR_188 ( );
FILL FILL_33_DFFSR_188 ( );
FILL FILL_34_DFFSR_188 ( );
FILL FILL_35_DFFSR_188 ( );
FILL FILL_36_DFFSR_188 ( );
FILL FILL_37_DFFSR_188 ( );
FILL FILL_38_DFFSR_188 ( );
FILL FILL_39_DFFSR_188 ( );
FILL FILL_40_DFFSR_188 ( );
FILL FILL_41_DFFSR_188 ( );
FILL FILL_42_DFFSR_188 ( );
FILL FILL_43_DFFSR_188 ( );
FILL FILL_44_DFFSR_188 ( );
FILL FILL_45_DFFSR_188 ( );
FILL FILL_46_DFFSR_188 ( );
FILL FILL_47_DFFSR_188 ( );
FILL FILL_48_DFFSR_188 ( );
FILL FILL_49_DFFSR_188 ( );
FILL FILL_50_DFFSR_188 ( );
FILL FILL_51_DFFSR_188 ( );
FILL FILL_0_DFFSR_203 ( );
FILL FILL_1_DFFSR_203 ( );
FILL FILL_2_DFFSR_203 ( );
FILL FILL_3_DFFSR_203 ( );
FILL FILL_4_DFFSR_203 ( );
FILL FILL_5_DFFSR_203 ( );
FILL FILL_6_DFFSR_203 ( );
FILL FILL_7_DFFSR_203 ( );
FILL FILL_8_DFFSR_203 ( );
FILL FILL_9_DFFSR_203 ( );
FILL FILL_10_DFFSR_203 ( );
FILL FILL_11_DFFSR_203 ( );
FILL FILL_12_DFFSR_203 ( );
FILL FILL_13_DFFSR_203 ( );
FILL FILL_14_DFFSR_203 ( );
FILL FILL_15_DFFSR_203 ( );
FILL FILL_16_DFFSR_203 ( );
FILL FILL_17_DFFSR_203 ( );
FILL FILL_18_DFFSR_203 ( );
FILL FILL_19_DFFSR_203 ( );
FILL FILL_20_DFFSR_203 ( );
FILL FILL_21_DFFSR_203 ( );
FILL FILL_22_DFFSR_203 ( );
FILL FILL_23_DFFSR_203 ( );
FILL FILL_24_DFFSR_203 ( );
FILL FILL_25_DFFSR_203 ( );
FILL FILL_26_DFFSR_203 ( );
FILL FILL_27_DFFSR_203 ( );
FILL FILL_28_DFFSR_203 ( );
FILL FILL_29_DFFSR_203 ( );
FILL FILL_30_DFFSR_203 ( );
FILL FILL_31_DFFSR_203 ( );
FILL FILL_32_DFFSR_203 ( );
FILL FILL_33_DFFSR_203 ( );
FILL FILL_34_DFFSR_203 ( );
FILL FILL_35_DFFSR_203 ( );
FILL FILL_36_DFFSR_203 ( );
FILL FILL_37_DFFSR_203 ( );
FILL FILL_38_DFFSR_203 ( );
FILL FILL_39_DFFSR_203 ( );
FILL FILL_40_DFFSR_203 ( );
FILL FILL_41_DFFSR_203 ( );
FILL FILL_42_DFFSR_203 ( );
FILL FILL_43_DFFSR_203 ( );
FILL FILL_44_DFFSR_203 ( );
FILL FILL_45_DFFSR_203 ( );
FILL FILL_46_DFFSR_203 ( );
FILL FILL_47_DFFSR_203 ( );
FILL FILL_48_DFFSR_203 ( );
FILL FILL_49_DFFSR_203 ( );
FILL FILL_50_DFFSR_203 ( );
FILL FILL_0_AND2X2_14 ( );
FILL FILL_1_AND2X2_14 ( );
FILL FILL_2_AND2X2_14 ( );
FILL FILL_3_AND2X2_14 ( );
FILL FILL_4_AND2X2_14 ( );
FILL FILL_5_AND2X2_14 ( );
FILL FILL_6_AND2X2_14 ( );
FILL FILL_7_AND2X2_14 ( );
FILL FILL_8_AND2X2_14 ( );
FILL FILL_9_AND2X2_14 ( );
FILL FILL_0_BUFX2_34 ( );
FILL FILL_1_BUFX2_34 ( );
FILL FILL_2_BUFX2_34 ( );
FILL FILL_3_BUFX2_34 ( );
FILL FILL_4_BUFX2_34 ( );
FILL FILL_5_BUFX2_34 ( );
FILL FILL_6_BUFX2_34 ( );
FILL FILL_0_DFFSR_177 ( );
FILL FILL_1_DFFSR_177 ( );
FILL FILL_2_DFFSR_177 ( );
FILL FILL_3_DFFSR_177 ( );
FILL FILL_4_DFFSR_177 ( );
FILL FILL_5_DFFSR_177 ( );
FILL FILL_6_DFFSR_177 ( );
FILL FILL_7_DFFSR_177 ( );
FILL FILL_8_DFFSR_177 ( );
FILL FILL_9_DFFSR_177 ( );
FILL FILL_10_DFFSR_177 ( );
FILL FILL_11_DFFSR_177 ( );
FILL FILL_12_DFFSR_177 ( );
FILL FILL_13_DFFSR_177 ( );
FILL FILL_14_DFFSR_177 ( );
FILL FILL_15_DFFSR_177 ( );
FILL FILL_16_DFFSR_177 ( );
FILL FILL_17_DFFSR_177 ( );
FILL FILL_18_DFFSR_177 ( );
FILL FILL_19_DFFSR_177 ( );
FILL FILL_20_DFFSR_177 ( );
FILL FILL_21_DFFSR_177 ( );
FILL FILL_22_DFFSR_177 ( );
FILL FILL_23_DFFSR_177 ( );
FILL FILL_24_DFFSR_177 ( );
FILL FILL_25_DFFSR_177 ( );
FILL FILL_26_DFFSR_177 ( );
FILL FILL_27_DFFSR_177 ( );
FILL FILL_28_DFFSR_177 ( );
FILL FILL_29_DFFSR_177 ( );
FILL FILL_30_DFFSR_177 ( );
FILL FILL_31_DFFSR_177 ( );
FILL FILL_32_DFFSR_177 ( );
FILL FILL_33_DFFSR_177 ( );
FILL FILL_34_DFFSR_177 ( );
FILL FILL_35_DFFSR_177 ( );
FILL FILL_36_DFFSR_177 ( );
FILL FILL_37_DFFSR_177 ( );
FILL FILL_38_DFFSR_177 ( );
FILL FILL_39_DFFSR_177 ( );
FILL FILL_40_DFFSR_177 ( );
FILL FILL_41_DFFSR_177 ( );
FILL FILL_42_DFFSR_177 ( );
FILL FILL_43_DFFSR_177 ( );
FILL FILL_44_DFFSR_177 ( );
FILL FILL_45_DFFSR_177 ( );
FILL FILL_46_DFFSR_177 ( );
FILL FILL_47_DFFSR_177 ( );
FILL FILL_48_DFFSR_177 ( );
FILL FILL_49_DFFSR_177 ( );
FILL FILL_50_DFFSR_177 ( );
FILL FILL_0_BUFX2_31 ( );
FILL FILL_1_BUFX2_31 ( );
FILL FILL_2_BUFX2_31 ( );
FILL FILL_3_BUFX2_31 ( );
FILL FILL_4_BUFX2_31 ( );
FILL FILL_5_BUFX2_31 ( );
FILL FILL_6_BUFX2_31 ( );
FILL FILL_0_AOI22X1_15 ( );
FILL FILL_1_AOI22X1_15 ( );
FILL FILL_2_AOI22X1_15 ( );
FILL FILL_3_AOI22X1_15 ( );
FILL FILL_4_AOI22X1_15 ( );
FILL FILL_5_AOI22X1_15 ( );
FILL FILL_6_AOI22X1_15 ( );
FILL FILL_7_AOI22X1_15 ( );
FILL FILL_8_AOI22X1_15 ( );
FILL FILL_9_AOI22X1_15 ( );
FILL FILL_10_AOI22X1_15 ( );
FILL FILL_11_AOI22X1_15 ( );
FILL FILL_0_NAND3X1_119 ( );
FILL FILL_1_NAND3X1_119 ( );
FILL FILL_2_NAND3X1_119 ( );
FILL FILL_3_NAND3X1_119 ( );
FILL FILL_4_NAND3X1_119 ( );
FILL FILL_5_NAND3X1_119 ( );
FILL FILL_6_NAND3X1_119 ( );
FILL FILL_7_NAND3X1_119 ( );
FILL FILL_8_NAND3X1_119 ( );
FILL FILL_0_NAND3X1_116 ( );
FILL FILL_1_NAND3X1_116 ( );
FILL FILL_2_NAND3X1_116 ( );
FILL FILL_3_NAND3X1_116 ( );
FILL FILL_4_NAND3X1_116 ( );
FILL FILL_5_NAND3X1_116 ( );
FILL FILL_6_NAND3X1_116 ( );
FILL FILL_7_NAND3X1_116 ( );
FILL FILL_8_NAND3X1_116 ( );
FILL FILL_0_DFFSR_232 ( );
FILL FILL_1_DFFSR_232 ( );
FILL FILL_2_DFFSR_232 ( );
FILL FILL_3_DFFSR_232 ( );
FILL FILL_4_DFFSR_232 ( );
FILL FILL_5_DFFSR_232 ( );
FILL FILL_6_DFFSR_232 ( );
FILL FILL_7_DFFSR_232 ( );
FILL FILL_8_DFFSR_232 ( );
FILL FILL_9_DFFSR_232 ( );
FILL FILL_10_DFFSR_232 ( );
FILL FILL_11_DFFSR_232 ( );
FILL FILL_12_DFFSR_232 ( );
FILL FILL_13_DFFSR_232 ( );
FILL FILL_14_DFFSR_232 ( );
FILL FILL_15_DFFSR_232 ( );
FILL FILL_16_DFFSR_232 ( );
FILL FILL_17_DFFSR_232 ( );
FILL FILL_18_DFFSR_232 ( );
FILL FILL_19_DFFSR_232 ( );
FILL FILL_20_DFFSR_232 ( );
FILL FILL_21_DFFSR_232 ( );
FILL FILL_22_DFFSR_232 ( );
FILL FILL_23_DFFSR_232 ( );
FILL FILL_24_DFFSR_232 ( );
FILL FILL_25_DFFSR_232 ( );
FILL FILL_26_DFFSR_232 ( );
FILL FILL_27_DFFSR_232 ( );
FILL FILL_28_DFFSR_232 ( );
FILL FILL_29_DFFSR_232 ( );
FILL FILL_30_DFFSR_232 ( );
FILL FILL_31_DFFSR_232 ( );
FILL FILL_32_DFFSR_232 ( );
FILL FILL_33_DFFSR_232 ( );
FILL FILL_34_DFFSR_232 ( );
FILL FILL_35_DFFSR_232 ( );
FILL FILL_36_DFFSR_232 ( );
FILL FILL_37_DFFSR_232 ( );
FILL FILL_38_DFFSR_232 ( );
FILL FILL_39_DFFSR_232 ( );
FILL FILL_40_DFFSR_232 ( );
FILL FILL_41_DFFSR_232 ( );
FILL FILL_42_DFFSR_232 ( );
FILL FILL_43_DFFSR_232 ( );
FILL FILL_44_DFFSR_232 ( );
FILL FILL_45_DFFSR_232 ( );
FILL FILL_46_DFFSR_232 ( );
FILL FILL_47_DFFSR_232 ( );
FILL FILL_48_DFFSR_232 ( );
FILL FILL_49_DFFSR_232 ( );
FILL FILL_50_DFFSR_232 ( );
FILL FILL_51_DFFSR_232 ( );
FILL FILL_0_NAND2X1_120 ( );
FILL FILL_1_NAND2X1_120 ( );
FILL FILL_2_NAND2X1_120 ( );
FILL FILL_3_NAND2X1_120 ( );
FILL FILL_4_NAND2X1_120 ( );
FILL FILL_5_NAND2X1_120 ( );
FILL FILL_6_NAND2X1_120 ( );
FILL FILL_0_NAND3X1_181 ( );
FILL FILL_1_NAND3X1_181 ( );
FILL FILL_2_NAND3X1_181 ( );
FILL FILL_3_NAND3X1_181 ( );
FILL FILL_4_NAND3X1_181 ( );
FILL FILL_5_NAND3X1_181 ( );
FILL FILL_6_NAND3X1_181 ( );
FILL FILL_7_NAND3X1_181 ( );
FILL FILL_8_NAND3X1_181 ( );
FILL FILL_0_AOI21X1_21 ( );
FILL FILL_1_AOI21X1_21 ( );
FILL FILL_2_AOI21X1_21 ( );
FILL FILL_3_AOI21X1_21 ( );
FILL FILL_4_AOI21X1_21 ( );
FILL FILL_5_AOI21X1_21 ( );
FILL FILL_6_AOI21X1_21 ( );
FILL FILL_7_AOI21X1_21 ( );
FILL FILL_8_AOI21X1_21 ( );
FILL FILL_0_OAI21X1_58 ( );
FILL FILL_1_OAI21X1_58 ( );
FILL FILL_2_OAI21X1_58 ( );
FILL FILL_3_OAI21X1_58 ( );
FILL FILL_4_OAI21X1_58 ( );
FILL FILL_5_OAI21X1_58 ( );
FILL FILL_6_OAI21X1_58 ( );
FILL FILL_7_OAI21X1_58 ( );
FILL FILL_8_OAI21X1_58 ( );
FILL FILL_9_OAI21X1_58 ( );
FILL FILL_0_NAND3X1_212 ( );
FILL FILL_1_NAND3X1_212 ( );
FILL FILL_2_NAND3X1_212 ( );
FILL FILL_3_NAND3X1_212 ( );
FILL FILL_4_NAND3X1_212 ( );
FILL FILL_5_NAND3X1_212 ( );
FILL FILL_6_NAND3X1_212 ( );
FILL FILL_7_NAND3X1_212 ( );
FILL FILL_8_NAND3X1_212 ( );
FILL FILL_0_NAND2X1_101 ( );
FILL FILL_1_NAND2X1_101 ( );
FILL FILL_2_NAND2X1_101 ( );
FILL FILL_3_NAND2X1_101 ( );
FILL FILL_4_NAND2X1_101 ( );
FILL FILL_5_NAND2X1_101 ( );
FILL FILL_6_NAND2X1_101 ( );
FILL FILL_0_NAND3X1_213 ( );
FILL FILL_1_NAND3X1_213 ( );
FILL FILL_2_NAND3X1_213 ( );
FILL FILL_3_NAND3X1_213 ( );
FILL FILL_4_NAND3X1_213 ( );
FILL FILL_5_NAND3X1_213 ( );
FILL FILL_6_NAND3X1_213 ( );
FILL FILL_7_NAND3X1_213 ( );
FILL FILL_8_NAND3X1_213 ( );
FILL FILL_0_AOI21X1_40 ( );
FILL FILL_1_AOI21X1_40 ( );
FILL FILL_2_AOI21X1_40 ( );
FILL FILL_3_AOI21X1_40 ( );
FILL FILL_4_AOI21X1_40 ( );
FILL FILL_5_AOI21X1_40 ( );
FILL FILL_6_AOI21X1_40 ( );
FILL FILL_7_AOI21X1_40 ( );
FILL FILL_8_AOI21X1_40 ( );
FILL FILL_9_AOI21X1_40 ( );
FILL FILL_0_NAND3X1_224 ( );
FILL FILL_1_NAND3X1_224 ( );
FILL FILL_2_NAND3X1_224 ( );
FILL FILL_3_NAND3X1_224 ( );
FILL FILL_4_NAND3X1_224 ( );
FILL FILL_5_NAND3X1_224 ( );
FILL FILL_6_NAND3X1_224 ( );
FILL FILL_7_NAND3X1_224 ( );
FILL FILL_8_NAND3X1_224 ( );
FILL FILL_0_NAND2X1_99 ( );
FILL FILL_1_NAND2X1_99 ( );
FILL FILL_2_NAND2X1_99 ( );
FILL FILL_3_NAND2X1_99 ( );
FILL FILL_4_NAND2X1_99 ( );
FILL FILL_5_NAND2X1_99 ( );
FILL FILL_6_NAND2X1_99 ( );
FILL FILL_0_OAI22X1_51 ( );
FILL FILL_1_OAI22X1_51 ( );
FILL FILL_2_OAI22X1_51 ( );
FILL FILL_3_OAI22X1_51 ( );
FILL FILL_4_OAI22X1_51 ( );
FILL FILL_5_OAI22X1_51 ( );
FILL FILL_6_OAI22X1_51 ( );
FILL FILL_7_OAI22X1_51 ( );
FILL FILL_8_OAI22X1_51 ( );
FILL FILL_9_OAI22X1_51 ( );
FILL FILL_10_OAI22X1_51 ( );
FILL FILL_11_OAI22X1_51 ( );
FILL FILL_0_NAND2X1_100 ( );
FILL FILL_1_NAND2X1_100 ( );
FILL FILL_2_NAND2X1_100 ( );
FILL FILL_3_NAND2X1_100 ( );
FILL FILL_4_NAND2X1_100 ( );
FILL FILL_5_NAND2X1_100 ( );
FILL FILL_6_NAND2X1_100 ( );
FILL FILL_0_OAI21X1_75 ( );
FILL FILL_1_OAI21X1_75 ( );
FILL FILL_2_OAI21X1_75 ( );
FILL FILL_3_OAI21X1_75 ( );
FILL FILL_4_OAI21X1_75 ( );
FILL FILL_5_OAI21X1_75 ( );
FILL FILL_6_OAI21X1_75 ( );
FILL FILL_7_OAI21X1_75 ( );
FILL FILL_8_OAI21X1_75 ( );
FILL FILL_0_INVX1_163 ( );
FILL FILL_1_INVX1_163 ( );
FILL FILL_2_INVX1_163 ( );
FILL FILL_3_INVX1_163 ( );
FILL FILL_0_AOI21X1_35 ( );
FILL FILL_1_AOI21X1_35 ( );
FILL FILL_2_AOI21X1_35 ( );
FILL FILL_3_AOI21X1_35 ( );
FILL FILL_4_AOI21X1_35 ( );
FILL FILL_5_AOI21X1_35 ( );
FILL FILL_6_AOI21X1_35 ( );
FILL FILL_7_AOI21X1_35 ( );
FILL FILL_8_AOI21X1_35 ( );
FILL FILL_9_AOI21X1_35 ( );
FILL FILL_0_NAND2X1_91 ( );
FILL FILL_1_NAND2X1_91 ( );
FILL FILL_2_NAND2X1_91 ( );
FILL FILL_3_NAND2X1_91 ( );
FILL FILL_4_NAND2X1_91 ( );
FILL FILL_5_NAND2X1_91 ( );
FILL FILL_6_NAND2X1_91 ( );
FILL FILL_0_DFFSR_270 ( );
FILL FILL_1_DFFSR_270 ( );
FILL FILL_2_DFFSR_270 ( );
FILL FILL_3_DFFSR_270 ( );
FILL FILL_4_DFFSR_270 ( );
FILL FILL_5_DFFSR_270 ( );
FILL FILL_6_DFFSR_270 ( );
FILL FILL_7_DFFSR_270 ( );
FILL FILL_8_DFFSR_270 ( );
FILL FILL_9_DFFSR_270 ( );
FILL FILL_10_DFFSR_270 ( );
FILL FILL_11_DFFSR_270 ( );
FILL FILL_12_DFFSR_270 ( );
FILL FILL_13_DFFSR_270 ( );
FILL FILL_14_DFFSR_270 ( );
FILL FILL_15_DFFSR_270 ( );
FILL FILL_16_DFFSR_270 ( );
FILL FILL_17_DFFSR_270 ( );
FILL FILL_18_DFFSR_270 ( );
FILL FILL_19_DFFSR_270 ( );
FILL FILL_20_DFFSR_270 ( );
FILL FILL_21_DFFSR_270 ( );
FILL FILL_22_DFFSR_270 ( );
FILL FILL_23_DFFSR_270 ( );
FILL FILL_24_DFFSR_270 ( );
FILL FILL_25_DFFSR_270 ( );
FILL FILL_26_DFFSR_270 ( );
FILL FILL_27_DFFSR_270 ( );
FILL FILL_28_DFFSR_270 ( );
FILL FILL_29_DFFSR_270 ( );
FILL FILL_30_DFFSR_270 ( );
FILL FILL_31_DFFSR_270 ( );
FILL FILL_32_DFFSR_270 ( );
FILL FILL_33_DFFSR_270 ( );
FILL FILL_34_DFFSR_270 ( );
FILL FILL_35_DFFSR_270 ( );
FILL FILL_36_DFFSR_270 ( );
FILL FILL_37_DFFSR_270 ( );
FILL FILL_38_DFFSR_270 ( );
FILL FILL_39_DFFSR_270 ( );
FILL FILL_40_DFFSR_270 ( );
FILL FILL_41_DFFSR_270 ( );
FILL FILL_42_DFFSR_270 ( );
FILL FILL_43_DFFSR_270 ( );
FILL FILL_44_DFFSR_270 ( );
FILL FILL_45_DFFSR_270 ( );
FILL FILL_46_DFFSR_270 ( );
FILL FILL_47_DFFSR_270 ( );
FILL FILL_48_DFFSR_270 ( );
FILL FILL_49_DFFSR_270 ( );
FILL FILL_50_DFFSR_270 ( );
FILL FILL_0_DFFPOSX1_35 ( );
FILL FILL_1_DFFPOSX1_35 ( );
FILL FILL_2_DFFPOSX1_35 ( );
FILL FILL_3_DFFPOSX1_35 ( );
FILL FILL_4_DFFPOSX1_35 ( );
FILL FILL_5_DFFPOSX1_35 ( );
FILL FILL_6_DFFPOSX1_35 ( );
FILL FILL_7_DFFPOSX1_35 ( );
FILL FILL_8_DFFPOSX1_35 ( );
FILL FILL_9_DFFPOSX1_35 ( );
FILL FILL_10_DFFPOSX1_35 ( );
FILL FILL_11_DFFPOSX1_35 ( );
FILL FILL_12_DFFPOSX1_35 ( );
FILL FILL_13_DFFPOSX1_35 ( );
FILL FILL_14_DFFPOSX1_35 ( );
FILL FILL_15_DFFPOSX1_35 ( );
FILL FILL_16_DFFPOSX1_35 ( );
FILL FILL_17_DFFPOSX1_35 ( );
FILL FILL_18_DFFPOSX1_35 ( );
FILL FILL_19_DFFPOSX1_35 ( );
FILL FILL_20_DFFPOSX1_35 ( );
FILL FILL_21_DFFPOSX1_35 ( );
FILL FILL_22_DFFPOSX1_35 ( );
FILL FILL_23_DFFPOSX1_35 ( );
FILL FILL_24_DFFPOSX1_35 ( );
FILL FILL_25_DFFPOSX1_35 ( );
FILL FILL_26_DFFPOSX1_35 ( );
FILL FILL_27_DFFPOSX1_35 ( );
FILL FILL_0_DFFSR_54 ( );
FILL FILL_1_DFFSR_54 ( );
FILL FILL_2_DFFSR_54 ( );
FILL FILL_3_DFFSR_54 ( );
FILL FILL_4_DFFSR_54 ( );
FILL FILL_5_DFFSR_54 ( );
FILL FILL_6_DFFSR_54 ( );
FILL FILL_7_DFFSR_54 ( );
FILL FILL_8_DFFSR_54 ( );
FILL FILL_9_DFFSR_54 ( );
FILL FILL_10_DFFSR_54 ( );
FILL FILL_11_DFFSR_54 ( );
FILL FILL_12_DFFSR_54 ( );
FILL FILL_13_DFFSR_54 ( );
FILL FILL_14_DFFSR_54 ( );
FILL FILL_15_DFFSR_54 ( );
FILL FILL_16_DFFSR_54 ( );
FILL FILL_17_DFFSR_54 ( );
FILL FILL_18_DFFSR_54 ( );
FILL FILL_19_DFFSR_54 ( );
FILL FILL_20_DFFSR_54 ( );
FILL FILL_21_DFFSR_54 ( );
FILL FILL_22_DFFSR_54 ( );
FILL FILL_23_DFFSR_54 ( );
FILL FILL_24_DFFSR_54 ( );
FILL FILL_25_DFFSR_54 ( );
FILL FILL_26_DFFSR_54 ( );
FILL FILL_27_DFFSR_54 ( );
FILL FILL_28_DFFSR_54 ( );
FILL FILL_29_DFFSR_54 ( );
FILL FILL_30_DFFSR_54 ( );
FILL FILL_31_DFFSR_54 ( );
FILL FILL_32_DFFSR_54 ( );
FILL FILL_33_DFFSR_54 ( );
FILL FILL_34_DFFSR_54 ( );
FILL FILL_35_DFFSR_54 ( );
FILL FILL_36_DFFSR_54 ( );
FILL FILL_37_DFFSR_54 ( );
FILL FILL_38_DFFSR_54 ( );
FILL FILL_39_DFFSR_54 ( );
FILL FILL_40_DFFSR_54 ( );
FILL FILL_41_DFFSR_54 ( );
FILL FILL_42_DFFSR_54 ( );
FILL FILL_43_DFFSR_54 ( );
FILL FILL_44_DFFSR_54 ( );
FILL FILL_45_DFFSR_54 ( );
FILL FILL_46_DFFSR_54 ( );
FILL FILL_47_DFFSR_54 ( );
FILL FILL_48_DFFSR_54 ( );
FILL FILL_49_DFFSR_54 ( );
FILL FILL_50_DFFSR_54 ( );
FILL FILL_51_DFFSR_54 ( );
FILL FILL_0_OAI21X1_85 ( );
FILL FILL_1_OAI21X1_85 ( );
FILL FILL_2_OAI21X1_85 ( );
FILL FILL_3_OAI21X1_85 ( );
FILL FILL_4_OAI21X1_85 ( );
FILL FILL_5_OAI21X1_85 ( );
FILL FILL_6_OAI21X1_85 ( );
FILL FILL_7_OAI21X1_85 ( );
FILL FILL_8_OAI21X1_85 ( );
FILL FILL_0_OAI22X1_41 ( );
FILL FILL_1_OAI22X1_41 ( );
FILL FILL_2_OAI22X1_41 ( );
FILL FILL_3_OAI22X1_41 ( );
FILL FILL_4_OAI22X1_41 ( );
FILL FILL_5_OAI22X1_41 ( );
FILL FILL_6_OAI22X1_41 ( );
FILL FILL_7_OAI22X1_41 ( );
FILL FILL_8_OAI22X1_41 ( );
FILL FILL_9_OAI22X1_41 ( );
FILL FILL_10_OAI22X1_41 ( );
FILL FILL_11_OAI22X1_41 ( );
FILL FILL_0_INVX1_83 ( );
FILL FILL_1_INVX1_83 ( );
FILL FILL_2_INVX1_83 ( );
FILL FILL_3_INVX1_83 ( );
FILL FILL_0_NAND3X1_134 ( );
FILL FILL_1_NAND3X1_134 ( );
FILL FILL_2_NAND3X1_134 ( );
FILL FILL_3_NAND3X1_134 ( );
FILL FILL_4_NAND3X1_134 ( );
FILL FILL_5_NAND3X1_134 ( );
FILL FILL_6_NAND3X1_134 ( );
FILL FILL_7_NAND3X1_134 ( );
FILL FILL_8_NAND3X1_134 ( );
FILL FILL_0_INVX1_79 ( );
FILL FILL_1_INVX1_79 ( );
FILL FILL_2_INVX1_79 ( );
FILL FILL_3_INVX1_79 ( );
FILL FILL_0_OAI22X1_32 ( );
FILL FILL_1_OAI22X1_32 ( );
FILL FILL_2_OAI22X1_32 ( );
FILL FILL_3_OAI22X1_32 ( );
FILL FILL_4_OAI22X1_32 ( );
FILL FILL_5_OAI22X1_32 ( );
FILL FILL_6_OAI22X1_32 ( );
FILL FILL_7_OAI22X1_32 ( );
FILL FILL_8_OAI22X1_32 ( );
FILL FILL_9_OAI22X1_32 ( );
FILL FILL_10_OAI22X1_32 ( );
FILL FILL_11_OAI22X1_32 ( );
FILL FILL_0_NOR2X1_31 ( );
FILL FILL_1_NOR2X1_31 ( );
FILL FILL_2_NOR2X1_31 ( );
FILL FILL_3_NOR2X1_31 ( );
FILL FILL_4_NOR2X1_31 ( );
FILL FILL_5_NOR2X1_31 ( );
FILL FILL_6_NOR2X1_31 ( );
FILL FILL_0_DFFSR_185 ( );
FILL FILL_1_DFFSR_185 ( );
FILL FILL_2_DFFSR_185 ( );
FILL FILL_3_DFFSR_185 ( );
FILL FILL_4_DFFSR_185 ( );
FILL FILL_5_DFFSR_185 ( );
FILL FILL_6_DFFSR_185 ( );
FILL FILL_7_DFFSR_185 ( );
FILL FILL_8_DFFSR_185 ( );
FILL FILL_9_DFFSR_185 ( );
FILL FILL_10_DFFSR_185 ( );
FILL FILL_11_DFFSR_185 ( );
FILL FILL_12_DFFSR_185 ( );
FILL FILL_13_DFFSR_185 ( );
FILL FILL_14_DFFSR_185 ( );
FILL FILL_15_DFFSR_185 ( );
FILL FILL_16_DFFSR_185 ( );
FILL FILL_17_DFFSR_185 ( );
FILL FILL_18_DFFSR_185 ( );
FILL FILL_19_DFFSR_185 ( );
FILL FILL_20_DFFSR_185 ( );
FILL FILL_21_DFFSR_185 ( );
FILL FILL_22_DFFSR_185 ( );
FILL FILL_23_DFFSR_185 ( );
FILL FILL_24_DFFSR_185 ( );
FILL FILL_25_DFFSR_185 ( );
FILL FILL_26_DFFSR_185 ( );
FILL FILL_27_DFFSR_185 ( );
FILL FILL_28_DFFSR_185 ( );
FILL FILL_29_DFFSR_185 ( );
FILL FILL_30_DFFSR_185 ( );
FILL FILL_31_DFFSR_185 ( );
FILL FILL_32_DFFSR_185 ( );
FILL FILL_33_DFFSR_185 ( );
FILL FILL_34_DFFSR_185 ( );
FILL FILL_35_DFFSR_185 ( );
FILL FILL_36_DFFSR_185 ( );
FILL FILL_37_DFFSR_185 ( );
FILL FILL_38_DFFSR_185 ( );
FILL FILL_39_DFFSR_185 ( );
FILL FILL_40_DFFSR_185 ( );
FILL FILL_41_DFFSR_185 ( );
FILL FILL_42_DFFSR_185 ( );
FILL FILL_43_DFFSR_185 ( );
FILL FILL_44_DFFSR_185 ( );
FILL FILL_45_DFFSR_185 ( );
FILL FILL_46_DFFSR_185 ( );
FILL FILL_47_DFFSR_185 ( );
FILL FILL_48_DFFSR_185 ( );
FILL FILL_49_DFFSR_185 ( );
FILL FILL_50_DFFSR_185 ( );
FILL FILL_51_DFFSR_185 ( );
FILL FILL_0_INVX1_103 ( );
FILL FILL_1_INVX1_103 ( );
FILL FILL_2_INVX1_103 ( );
FILL FILL_3_INVX1_103 ( );
FILL FILL_4_INVX1_103 ( );
FILL FILL_0_INVX1_61 ( );
FILL FILL_1_INVX1_61 ( );
FILL FILL_2_INVX1_61 ( );
FILL FILL_3_INVX1_61 ( );
FILL FILL_4_INVX1_61 ( );
FILL FILL_0_OAI22X1_25 ( );
FILL FILL_1_OAI22X1_25 ( );
FILL FILL_2_OAI22X1_25 ( );
FILL FILL_3_OAI22X1_25 ( );
FILL FILL_4_OAI22X1_25 ( );
FILL FILL_5_OAI22X1_25 ( );
FILL FILL_6_OAI22X1_25 ( );
FILL FILL_7_OAI22X1_25 ( );
FILL FILL_8_OAI22X1_25 ( );
FILL FILL_9_OAI22X1_25 ( );
FILL FILL_10_OAI22X1_25 ( );
FILL FILL_0_AND2X2_25 ( );
FILL FILL_1_AND2X2_25 ( );
FILL FILL_2_AND2X2_25 ( );
FILL FILL_3_AND2X2_25 ( );
FILL FILL_4_AND2X2_25 ( );
FILL FILL_5_AND2X2_25 ( );
FILL FILL_6_AND2X2_25 ( );
FILL FILL_7_AND2X2_25 ( );
FILL FILL_8_AND2X2_25 ( );
FILL FILL_0_OAI22X1_26 ( );
FILL FILL_1_OAI22X1_26 ( );
FILL FILL_2_OAI22X1_26 ( );
FILL FILL_3_OAI22X1_26 ( );
FILL FILL_4_OAI22X1_26 ( );
FILL FILL_5_OAI22X1_26 ( );
FILL FILL_6_OAI22X1_26 ( );
FILL FILL_7_OAI22X1_26 ( );
FILL FILL_8_OAI22X1_26 ( );
FILL FILL_9_OAI22X1_26 ( );
FILL FILL_10_OAI22X1_26 ( );
FILL FILL_0_NOR2X1_55 ( );
FILL FILL_1_NOR2X1_55 ( );
FILL FILL_2_NOR2X1_55 ( );
FILL FILL_3_NOR2X1_55 ( );
FILL FILL_4_NOR2X1_55 ( );
FILL FILL_5_NOR2X1_55 ( );
FILL FILL_6_NOR2X1_55 ( );
FILL FILL_0_OAI21X1_13 ( );
FILL FILL_1_OAI21X1_13 ( );
FILL FILL_2_OAI21X1_13 ( );
FILL FILL_3_OAI21X1_13 ( );
FILL FILL_4_OAI21X1_13 ( );
FILL FILL_5_OAI21X1_13 ( );
FILL FILL_6_OAI21X1_13 ( );
FILL FILL_7_OAI21X1_13 ( );
FILL FILL_8_OAI21X1_13 ( );
FILL FILL_0_DFFSR_239 ( );
FILL FILL_1_DFFSR_239 ( );
FILL FILL_2_DFFSR_239 ( );
FILL FILL_3_DFFSR_239 ( );
FILL FILL_4_DFFSR_239 ( );
FILL FILL_5_DFFSR_239 ( );
FILL FILL_6_DFFSR_239 ( );
FILL FILL_7_DFFSR_239 ( );
FILL FILL_8_DFFSR_239 ( );
FILL FILL_9_DFFSR_239 ( );
FILL FILL_10_DFFSR_239 ( );
FILL FILL_11_DFFSR_239 ( );
FILL FILL_12_DFFSR_239 ( );
FILL FILL_13_DFFSR_239 ( );
FILL FILL_14_DFFSR_239 ( );
FILL FILL_15_DFFSR_239 ( );
FILL FILL_16_DFFSR_239 ( );
FILL FILL_17_DFFSR_239 ( );
FILL FILL_18_DFFSR_239 ( );
FILL FILL_19_DFFSR_239 ( );
FILL FILL_20_DFFSR_239 ( );
FILL FILL_21_DFFSR_239 ( );
FILL FILL_22_DFFSR_239 ( );
FILL FILL_23_DFFSR_239 ( );
FILL FILL_24_DFFSR_239 ( );
FILL FILL_25_DFFSR_239 ( );
FILL FILL_26_DFFSR_239 ( );
FILL FILL_27_DFFSR_239 ( );
FILL FILL_28_DFFSR_239 ( );
FILL FILL_29_DFFSR_239 ( );
FILL FILL_30_DFFSR_239 ( );
FILL FILL_31_DFFSR_239 ( );
FILL FILL_32_DFFSR_239 ( );
FILL FILL_33_DFFSR_239 ( );
FILL FILL_34_DFFSR_239 ( );
FILL FILL_35_DFFSR_239 ( );
FILL FILL_36_DFFSR_239 ( );
FILL FILL_37_DFFSR_239 ( );
FILL FILL_38_DFFSR_239 ( );
FILL FILL_39_DFFSR_239 ( );
FILL FILL_40_DFFSR_239 ( );
FILL FILL_41_DFFSR_239 ( );
FILL FILL_42_DFFSR_239 ( );
FILL FILL_43_DFFSR_239 ( );
FILL FILL_44_DFFSR_239 ( );
FILL FILL_45_DFFSR_239 ( );
FILL FILL_46_DFFSR_239 ( );
FILL FILL_47_DFFSR_239 ( );
FILL FILL_48_DFFSR_239 ( );
FILL FILL_49_DFFSR_239 ( );
FILL FILL_50_DFFSR_239 ( );
FILL FILL_51_DFFSR_239 ( );
FILL FILL_0_INVX1_158 ( );
FILL FILL_1_INVX1_158 ( );
FILL FILL_2_INVX1_158 ( );
FILL FILL_3_INVX1_158 ( );
FILL FILL_4_INVX1_158 ( );
FILL FILL_0_AOI22X1_23 ( );
FILL FILL_1_AOI22X1_23 ( );
FILL FILL_2_AOI22X1_23 ( );
FILL FILL_3_AOI22X1_23 ( );
FILL FILL_4_AOI22X1_23 ( );
FILL FILL_5_AOI22X1_23 ( );
FILL FILL_6_AOI22X1_23 ( );
FILL FILL_7_AOI22X1_23 ( );
FILL FILL_8_AOI22X1_23 ( );
FILL FILL_9_AOI22X1_23 ( );
FILL FILL_10_AOI22X1_23 ( );
FILL FILL_11_AOI22X1_23 ( );
FILL FILL_0_AOI21X1_31 ( );
FILL FILL_1_AOI21X1_31 ( );
FILL FILL_2_AOI21X1_31 ( );
FILL FILL_3_AOI21X1_31 ( );
FILL FILL_4_AOI21X1_31 ( );
FILL FILL_5_AOI21X1_31 ( );
FILL FILL_6_AOI21X1_31 ( );
FILL FILL_7_AOI21X1_31 ( );
FILL FILL_8_AOI21X1_31 ( );
FILL FILL_0_NAND3X1_165 ( );
FILL FILL_1_NAND3X1_165 ( );
FILL FILL_2_NAND3X1_165 ( );
FILL FILL_3_NAND3X1_165 ( );
FILL FILL_4_NAND3X1_165 ( );
FILL FILL_5_NAND3X1_165 ( );
FILL FILL_6_NAND3X1_165 ( );
FILL FILL_7_NAND3X1_165 ( );
FILL FILL_8_NAND3X1_165 ( );
FILL FILL_0_AOI22X1_20 ( );
FILL FILL_1_AOI22X1_20 ( );
FILL FILL_2_AOI22X1_20 ( );
FILL FILL_3_AOI22X1_20 ( );
FILL FILL_4_AOI22X1_20 ( );
FILL FILL_5_AOI22X1_20 ( );
FILL FILL_6_AOI22X1_20 ( );
FILL FILL_7_AOI22X1_20 ( );
FILL FILL_8_AOI22X1_20 ( );
FILL FILL_9_AOI22X1_20 ( );
FILL FILL_10_AOI22X1_20 ( );
FILL FILL_11_AOI22X1_20 ( );
FILL FILL_0_AOI21X1_41 ( );
FILL FILL_1_AOI21X1_41 ( );
FILL FILL_2_AOI21X1_41 ( );
FILL FILL_3_AOI21X1_41 ( );
FILL FILL_4_AOI21X1_41 ( );
FILL FILL_5_AOI21X1_41 ( );
FILL FILL_6_AOI21X1_41 ( );
FILL FILL_7_AOI21X1_41 ( );
FILL FILL_8_AOI21X1_41 ( );
FILL FILL_0_INVX1_169 ( );
FILL FILL_1_INVX1_169 ( );
FILL FILL_2_INVX1_169 ( );
FILL FILL_3_INVX1_169 ( );
FILL FILL_4_INVX1_169 ( );
FILL FILL_0_DFFPOSX1_42 ( );
FILL FILL_1_DFFPOSX1_42 ( );
FILL FILL_2_DFFPOSX1_42 ( );
FILL FILL_3_DFFPOSX1_42 ( );
FILL FILL_4_DFFPOSX1_42 ( );
FILL FILL_5_DFFPOSX1_42 ( );
FILL FILL_6_DFFPOSX1_42 ( );
FILL FILL_7_DFFPOSX1_42 ( );
FILL FILL_8_DFFPOSX1_42 ( );
FILL FILL_9_DFFPOSX1_42 ( );
FILL FILL_10_DFFPOSX1_42 ( );
FILL FILL_11_DFFPOSX1_42 ( );
FILL FILL_12_DFFPOSX1_42 ( );
FILL FILL_13_DFFPOSX1_42 ( );
FILL FILL_14_DFFPOSX1_42 ( );
FILL FILL_15_DFFPOSX1_42 ( );
FILL FILL_16_DFFPOSX1_42 ( );
FILL FILL_17_DFFPOSX1_42 ( );
FILL FILL_18_DFFPOSX1_42 ( );
FILL FILL_19_DFFPOSX1_42 ( );
FILL FILL_20_DFFPOSX1_42 ( );
FILL FILL_21_DFFPOSX1_42 ( );
FILL FILL_22_DFFPOSX1_42 ( );
FILL FILL_23_DFFPOSX1_42 ( );
FILL FILL_24_DFFPOSX1_42 ( );
FILL FILL_25_DFFPOSX1_42 ( );
FILL FILL_26_DFFPOSX1_42 ( );
FILL FILL_27_DFFPOSX1_42 ( );
FILL FILL_0_AOI21X1_34 ( );
FILL FILL_1_AOI21X1_34 ( );
FILL FILL_2_AOI21X1_34 ( );
FILL FILL_3_AOI21X1_34 ( );
FILL FILL_4_AOI21X1_34 ( );
FILL FILL_5_AOI21X1_34 ( );
FILL FILL_6_AOI21X1_34 ( );
FILL FILL_7_AOI21X1_34 ( );
FILL FILL_8_AOI21X1_34 ( );
FILL FILL_0_DFFPOSX1_46 ( );
FILL FILL_1_DFFPOSX1_46 ( );
FILL FILL_2_DFFPOSX1_46 ( );
FILL FILL_3_DFFPOSX1_46 ( );
FILL FILL_4_DFFPOSX1_46 ( );
FILL FILL_5_DFFPOSX1_46 ( );
FILL FILL_6_DFFPOSX1_46 ( );
FILL FILL_7_DFFPOSX1_46 ( );
FILL FILL_8_DFFPOSX1_46 ( );
FILL FILL_9_DFFPOSX1_46 ( );
FILL FILL_10_DFFPOSX1_46 ( );
FILL FILL_11_DFFPOSX1_46 ( );
FILL FILL_12_DFFPOSX1_46 ( );
FILL FILL_13_DFFPOSX1_46 ( );
FILL FILL_14_DFFPOSX1_46 ( );
FILL FILL_15_DFFPOSX1_46 ( );
FILL FILL_16_DFFPOSX1_46 ( );
FILL FILL_17_DFFPOSX1_46 ( );
FILL FILL_18_DFFPOSX1_46 ( );
FILL FILL_19_DFFPOSX1_46 ( );
FILL FILL_20_DFFPOSX1_46 ( );
FILL FILL_21_DFFPOSX1_46 ( );
FILL FILL_22_DFFPOSX1_46 ( );
FILL FILL_23_DFFPOSX1_46 ( );
FILL FILL_24_DFFPOSX1_46 ( );
FILL FILL_25_DFFPOSX1_46 ( );
FILL FILL_26_DFFPOSX1_46 ( );
FILL FILL_27_DFFPOSX1_46 ( );
FILL FILL_0_INVX1_162 ( );
FILL FILL_1_INVX1_162 ( );
FILL FILL_2_INVX1_162 ( );
FILL FILL_3_INVX1_162 ( );
FILL FILL_4_INVX1_162 ( );
FILL FILL_0_DFFPOSX1_3 ( );
FILL FILL_1_DFFPOSX1_3 ( );
FILL FILL_2_DFFPOSX1_3 ( );
FILL FILL_3_DFFPOSX1_3 ( );
FILL FILL_4_DFFPOSX1_3 ( );
FILL FILL_5_DFFPOSX1_3 ( );
FILL FILL_6_DFFPOSX1_3 ( );
FILL FILL_7_DFFPOSX1_3 ( );
FILL FILL_8_DFFPOSX1_3 ( );
FILL FILL_9_DFFPOSX1_3 ( );
FILL FILL_10_DFFPOSX1_3 ( );
FILL FILL_11_DFFPOSX1_3 ( );
FILL FILL_12_DFFPOSX1_3 ( );
FILL FILL_13_DFFPOSX1_3 ( );
FILL FILL_14_DFFPOSX1_3 ( );
FILL FILL_15_DFFPOSX1_3 ( );
FILL FILL_16_DFFPOSX1_3 ( );
FILL FILL_17_DFFPOSX1_3 ( );
FILL FILL_18_DFFPOSX1_3 ( );
FILL FILL_19_DFFPOSX1_3 ( );
FILL FILL_20_DFFPOSX1_3 ( );
FILL FILL_21_DFFPOSX1_3 ( );
FILL FILL_22_DFFPOSX1_3 ( );
FILL FILL_23_DFFPOSX1_3 ( );
FILL FILL_24_DFFPOSX1_3 ( );
FILL FILL_25_DFFPOSX1_3 ( );
FILL FILL_26_DFFPOSX1_3 ( );
FILL FILL_27_DFFPOSX1_3 ( );
FILL FILL_0_INVX1_208 ( );
FILL FILL_1_INVX1_208 ( );
FILL FILL_2_INVX1_208 ( );
FILL FILL_3_INVX1_208 ( );
FILL FILL_4_INVX1_208 ( );
FILL FILL_0_DFFPOSX1_1 ( );
FILL FILL_1_DFFPOSX1_1 ( );
FILL FILL_2_DFFPOSX1_1 ( );
FILL FILL_3_DFFPOSX1_1 ( );
FILL FILL_4_DFFPOSX1_1 ( );
FILL FILL_5_DFFPOSX1_1 ( );
FILL FILL_6_DFFPOSX1_1 ( );
FILL FILL_7_DFFPOSX1_1 ( );
FILL FILL_8_DFFPOSX1_1 ( );
FILL FILL_9_DFFPOSX1_1 ( );
FILL FILL_10_DFFPOSX1_1 ( );
FILL FILL_11_DFFPOSX1_1 ( );
FILL FILL_12_DFFPOSX1_1 ( );
FILL FILL_13_DFFPOSX1_1 ( );
FILL FILL_14_DFFPOSX1_1 ( );
FILL FILL_15_DFFPOSX1_1 ( );
FILL FILL_16_DFFPOSX1_1 ( );
FILL FILL_17_DFFPOSX1_1 ( );
FILL FILL_18_DFFPOSX1_1 ( );
FILL FILL_19_DFFPOSX1_1 ( );
FILL FILL_20_DFFPOSX1_1 ( );
FILL FILL_21_DFFPOSX1_1 ( );
FILL FILL_22_DFFPOSX1_1 ( );
FILL FILL_23_DFFPOSX1_1 ( );
FILL FILL_24_DFFPOSX1_1 ( );
FILL FILL_25_DFFPOSX1_1 ( );
FILL FILL_26_DFFPOSX1_1 ( );
FILL FILL_27_DFFPOSX1_1 ( );
FILL FILL_0_OAI21X1_18 ( );
FILL FILL_1_OAI21X1_18 ( );
FILL FILL_2_OAI21X1_18 ( );
FILL FILL_3_OAI21X1_18 ( );
FILL FILL_4_OAI21X1_18 ( );
FILL FILL_5_OAI21X1_18 ( );
FILL FILL_6_OAI21X1_18 ( );
FILL FILL_7_OAI21X1_18 ( );
FILL FILL_8_OAI21X1_18 ( );
FILL FILL_0_INVX1_39 ( );
FILL FILL_1_INVX1_39 ( );
FILL FILL_2_INVX1_39 ( );
FILL FILL_3_INVX1_39 ( );
FILL FILL_0_NOR2X1_77 ( );
FILL FILL_1_NOR2X1_77 ( );
FILL FILL_2_NOR2X1_77 ( );
FILL FILL_3_NOR2X1_77 ( );
FILL FILL_4_NOR2X1_77 ( );
FILL FILL_5_NOR2X1_77 ( );
FILL FILL_6_NOR2X1_77 ( );
FILL FILL_0_DFFSR_257 ( );
FILL FILL_1_DFFSR_257 ( );
FILL FILL_2_DFFSR_257 ( );
FILL FILL_3_DFFSR_257 ( );
FILL FILL_4_DFFSR_257 ( );
FILL FILL_5_DFFSR_257 ( );
FILL FILL_6_DFFSR_257 ( );
FILL FILL_7_DFFSR_257 ( );
FILL FILL_8_DFFSR_257 ( );
FILL FILL_9_DFFSR_257 ( );
FILL FILL_10_DFFSR_257 ( );
FILL FILL_11_DFFSR_257 ( );
FILL FILL_12_DFFSR_257 ( );
FILL FILL_13_DFFSR_257 ( );
FILL FILL_14_DFFSR_257 ( );
FILL FILL_15_DFFSR_257 ( );
FILL FILL_16_DFFSR_257 ( );
FILL FILL_17_DFFSR_257 ( );
FILL FILL_18_DFFSR_257 ( );
FILL FILL_19_DFFSR_257 ( );
FILL FILL_20_DFFSR_257 ( );
FILL FILL_21_DFFSR_257 ( );
FILL FILL_22_DFFSR_257 ( );
FILL FILL_23_DFFSR_257 ( );
FILL FILL_24_DFFSR_257 ( );
FILL FILL_25_DFFSR_257 ( );
FILL FILL_26_DFFSR_257 ( );
FILL FILL_27_DFFSR_257 ( );
FILL FILL_28_DFFSR_257 ( );
FILL FILL_29_DFFSR_257 ( );
FILL FILL_30_DFFSR_257 ( );
FILL FILL_31_DFFSR_257 ( );
FILL FILL_32_DFFSR_257 ( );
FILL FILL_33_DFFSR_257 ( );
FILL FILL_34_DFFSR_257 ( );
FILL FILL_35_DFFSR_257 ( );
FILL FILL_36_DFFSR_257 ( );
FILL FILL_37_DFFSR_257 ( );
FILL FILL_38_DFFSR_257 ( );
FILL FILL_39_DFFSR_257 ( );
FILL FILL_40_DFFSR_257 ( );
FILL FILL_41_DFFSR_257 ( );
FILL FILL_42_DFFSR_257 ( );
FILL FILL_43_DFFSR_257 ( );
FILL FILL_44_DFFSR_257 ( );
FILL FILL_45_DFFSR_257 ( );
FILL FILL_46_DFFSR_257 ( );
FILL FILL_47_DFFSR_257 ( );
FILL FILL_48_DFFSR_257 ( );
FILL FILL_49_DFFSR_257 ( );
FILL FILL_50_DFFSR_257 ( );
FILL FILL_0_INVX1_84 ( );
FILL FILL_1_INVX1_84 ( );
FILL FILL_2_INVX1_84 ( );
FILL FILL_3_INVX1_84 ( );
FILL FILL_4_INVX1_84 ( );
FILL FILL_0_NOR2X1_50 ( );
FILL FILL_1_NOR2X1_50 ( );
FILL FILL_2_NOR2X1_50 ( );
FILL FILL_3_NOR2X1_50 ( );
FILL FILL_4_NOR2X1_50 ( );
FILL FILL_5_NOR2X1_50 ( );
FILL FILL_6_NOR2X1_50 ( );
FILL FILL_0_NAND2X1_44 ( );
FILL FILL_1_NAND2X1_44 ( );
FILL FILL_2_NAND2X1_44 ( );
FILL FILL_3_NAND2X1_44 ( );
FILL FILL_4_NAND2X1_44 ( );
FILL FILL_5_NAND2X1_44 ( );
FILL FILL_6_NAND2X1_44 ( );
FILL FILL_0_NAND2X1_55 ( );
FILL FILL_1_NAND2X1_55 ( );
FILL FILL_2_NAND2X1_55 ( );
FILL FILL_3_NAND2X1_55 ( );
FILL FILL_4_NAND2X1_55 ( );
FILL FILL_5_NAND2X1_55 ( );
FILL FILL_6_NAND2X1_55 ( );
FILL FILL_0_DFFSR_190 ( );
FILL FILL_1_DFFSR_190 ( );
FILL FILL_2_DFFSR_190 ( );
FILL FILL_3_DFFSR_190 ( );
FILL FILL_4_DFFSR_190 ( );
FILL FILL_5_DFFSR_190 ( );
FILL FILL_6_DFFSR_190 ( );
FILL FILL_7_DFFSR_190 ( );
FILL FILL_8_DFFSR_190 ( );
FILL FILL_9_DFFSR_190 ( );
FILL FILL_10_DFFSR_190 ( );
FILL FILL_11_DFFSR_190 ( );
FILL FILL_12_DFFSR_190 ( );
FILL FILL_13_DFFSR_190 ( );
FILL FILL_14_DFFSR_190 ( );
FILL FILL_15_DFFSR_190 ( );
FILL FILL_16_DFFSR_190 ( );
FILL FILL_17_DFFSR_190 ( );
FILL FILL_18_DFFSR_190 ( );
FILL FILL_19_DFFSR_190 ( );
FILL FILL_20_DFFSR_190 ( );
FILL FILL_21_DFFSR_190 ( );
FILL FILL_22_DFFSR_190 ( );
FILL FILL_23_DFFSR_190 ( );
FILL FILL_24_DFFSR_190 ( );
FILL FILL_25_DFFSR_190 ( );
FILL FILL_26_DFFSR_190 ( );
FILL FILL_27_DFFSR_190 ( );
FILL FILL_28_DFFSR_190 ( );
FILL FILL_29_DFFSR_190 ( );
FILL FILL_30_DFFSR_190 ( );
FILL FILL_31_DFFSR_190 ( );
FILL FILL_32_DFFSR_190 ( );
FILL FILL_33_DFFSR_190 ( );
FILL FILL_34_DFFSR_190 ( );
FILL FILL_35_DFFSR_190 ( );
FILL FILL_36_DFFSR_190 ( );
FILL FILL_37_DFFSR_190 ( );
FILL FILL_38_DFFSR_190 ( );
FILL FILL_39_DFFSR_190 ( );
FILL FILL_40_DFFSR_190 ( );
FILL FILL_41_DFFSR_190 ( );
FILL FILL_42_DFFSR_190 ( );
FILL FILL_43_DFFSR_190 ( );
FILL FILL_44_DFFSR_190 ( );
FILL FILL_45_DFFSR_190 ( );
FILL FILL_46_DFFSR_190 ( );
FILL FILL_47_DFFSR_190 ( );
FILL FILL_48_DFFSR_190 ( );
FILL FILL_49_DFFSR_190 ( );
FILL FILL_50_DFFSR_190 ( );
FILL FILL_0_NAND3X1_72 ( );
FILL FILL_1_NAND3X1_72 ( );
FILL FILL_2_NAND3X1_72 ( );
FILL FILL_3_NAND3X1_72 ( );
FILL FILL_4_NAND3X1_72 ( );
FILL FILL_5_NAND3X1_72 ( );
FILL FILL_6_NAND3X1_72 ( );
FILL FILL_7_NAND3X1_72 ( );
FILL FILL_8_NAND3X1_72 ( );
FILL FILL_0_INVX1_60 ( );
FILL FILL_1_INVX1_60 ( );
FILL FILL_2_INVX1_60 ( );
FILL FILL_3_INVX1_60 ( );
FILL FILL_4_INVX1_60 ( );
FILL FILL_0_DFFSR_223 ( );
FILL FILL_1_DFFSR_223 ( );
FILL FILL_2_DFFSR_223 ( );
FILL FILL_3_DFFSR_223 ( );
FILL FILL_4_DFFSR_223 ( );
FILL FILL_5_DFFSR_223 ( );
FILL FILL_6_DFFSR_223 ( );
FILL FILL_7_DFFSR_223 ( );
FILL FILL_8_DFFSR_223 ( );
FILL FILL_9_DFFSR_223 ( );
FILL FILL_10_DFFSR_223 ( );
FILL FILL_11_DFFSR_223 ( );
FILL FILL_12_DFFSR_223 ( );
FILL FILL_13_DFFSR_223 ( );
FILL FILL_14_DFFSR_223 ( );
FILL FILL_15_DFFSR_223 ( );
FILL FILL_16_DFFSR_223 ( );
FILL FILL_17_DFFSR_223 ( );
FILL FILL_18_DFFSR_223 ( );
FILL FILL_19_DFFSR_223 ( );
FILL FILL_20_DFFSR_223 ( );
FILL FILL_21_DFFSR_223 ( );
FILL FILL_22_DFFSR_223 ( );
FILL FILL_23_DFFSR_223 ( );
FILL FILL_24_DFFSR_223 ( );
FILL FILL_25_DFFSR_223 ( );
FILL FILL_26_DFFSR_223 ( );
FILL FILL_27_DFFSR_223 ( );
FILL FILL_28_DFFSR_223 ( );
FILL FILL_29_DFFSR_223 ( );
FILL FILL_30_DFFSR_223 ( );
FILL FILL_31_DFFSR_223 ( );
FILL FILL_32_DFFSR_223 ( );
FILL FILL_33_DFFSR_223 ( );
FILL FILL_34_DFFSR_223 ( );
FILL FILL_35_DFFSR_223 ( );
FILL FILL_36_DFFSR_223 ( );
FILL FILL_37_DFFSR_223 ( );
FILL FILL_38_DFFSR_223 ( );
FILL FILL_39_DFFSR_223 ( );
FILL FILL_40_DFFSR_223 ( );
FILL FILL_41_DFFSR_223 ( );
FILL FILL_42_DFFSR_223 ( );
FILL FILL_43_DFFSR_223 ( );
FILL FILL_44_DFFSR_223 ( );
FILL FILL_45_DFFSR_223 ( );
FILL FILL_46_DFFSR_223 ( );
FILL FILL_47_DFFSR_223 ( );
FILL FILL_48_DFFSR_223 ( );
FILL FILL_49_DFFSR_223 ( );
FILL FILL_50_DFFSR_223 ( );
FILL FILL_51_DFFSR_223 ( );
FILL FILL_0_NAND2X1_46 ( );
FILL FILL_1_NAND2X1_46 ( );
FILL FILL_2_NAND2X1_46 ( );
FILL FILL_3_NAND2X1_46 ( );
FILL FILL_4_NAND2X1_46 ( );
FILL FILL_5_NAND2X1_46 ( );
FILL FILL_6_NAND2X1_46 ( );
FILL FILL_0_NOR2X1_48 ( );
FILL FILL_1_NOR2X1_48 ( );
FILL FILL_2_NOR2X1_48 ( );
FILL FILL_3_NOR2X1_48 ( );
FILL FILL_4_NOR2X1_48 ( );
FILL FILL_5_NOR2X1_48 ( );
FILL FILL_6_NOR2X1_48 ( );
FILL FILL_0_NAND2X1_45 ( );
FILL FILL_1_NAND2X1_45 ( );
FILL FILL_2_NAND2X1_45 ( );
FILL FILL_3_NAND2X1_45 ( );
FILL FILL_4_NAND2X1_45 ( );
FILL FILL_5_NAND2X1_45 ( );
FILL FILL_6_NAND2X1_45 ( );
FILL FILL_0_DFFSR_240 ( );
FILL FILL_1_DFFSR_240 ( );
FILL FILL_2_DFFSR_240 ( );
FILL FILL_3_DFFSR_240 ( );
FILL FILL_4_DFFSR_240 ( );
FILL FILL_5_DFFSR_240 ( );
FILL FILL_6_DFFSR_240 ( );
FILL FILL_7_DFFSR_240 ( );
FILL FILL_8_DFFSR_240 ( );
FILL FILL_9_DFFSR_240 ( );
FILL FILL_10_DFFSR_240 ( );
FILL FILL_11_DFFSR_240 ( );
FILL FILL_12_DFFSR_240 ( );
FILL FILL_13_DFFSR_240 ( );
FILL FILL_14_DFFSR_240 ( );
FILL FILL_15_DFFSR_240 ( );
FILL FILL_16_DFFSR_240 ( );
FILL FILL_17_DFFSR_240 ( );
FILL FILL_18_DFFSR_240 ( );
FILL FILL_19_DFFSR_240 ( );
FILL FILL_20_DFFSR_240 ( );
FILL FILL_21_DFFSR_240 ( );
FILL FILL_22_DFFSR_240 ( );
FILL FILL_23_DFFSR_240 ( );
FILL FILL_24_DFFSR_240 ( );
FILL FILL_25_DFFSR_240 ( );
FILL FILL_26_DFFSR_240 ( );
FILL FILL_27_DFFSR_240 ( );
FILL FILL_28_DFFSR_240 ( );
FILL FILL_29_DFFSR_240 ( );
FILL FILL_30_DFFSR_240 ( );
FILL FILL_31_DFFSR_240 ( );
FILL FILL_32_DFFSR_240 ( );
FILL FILL_33_DFFSR_240 ( );
FILL FILL_34_DFFSR_240 ( );
FILL FILL_35_DFFSR_240 ( );
FILL FILL_36_DFFSR_240 ( );
FILL FILL_37_DFFSR_240 ( );
FILL FILL_38_DFFSR_240 ( );
FILL FILL_39_DFFSR_240 ( );
FILL FILL_40_DFFSR_240 ( );
FILL FILL_41_DFFSR_240 ( );
FILL FILL_42_DFFSR_240 ( );
FILL FILL_43_DFFSR_240 ( );
FILL FILL_44_DFFSR_240 ( );
FILL FILL_45_DFFSR_240 ( );
FILL FILL_46_DFFSR_240 ( );
FILL FILL_47_DFFSR_240 ( );
FILL FILL_48_DFFSR_240 ( );
FILL FILL_49_DFFSR_240 ( );
FILL FILL_50_DFFSR_240 ( );
FILL FILL_0_NAND3X1_171 ( );
FILL FILL_1_NAND3X1_171 ( );
FILL FILL_2_NAND3X1_171 ( );
FILL FILL_3_NAND3X1_171 ( );
FILL FILL_4_NAND3X1_171 ( );
FILL FILL_5_NAND3X1_171 ( );
FILL FILL_6_NAND3X1_171 ( );
FILL FILL_7_NAND3X1_171 ( );
FILL FILL_8_NAND3X1_171 ( );
FILL FILL_9_NAND3X1_171 ( );
FILL FILL_0_NAND2X1_83 ( );
FILL FILL_1_NAND2X1_83 ( );
FILL FILL_2_NAND2X1_83 ( );
FILL FILL_3_NAND2X1_83 ( );
FILL FILL_4_NAND2X1_83 ( );
FILL FILL_5_NAND2X1_83 ( );
FILL FILL_6_NAND2X1_83 ( );
FILL FILL_0_AND2X2_35 ( );
FILL FILL_1_AND2X2_35 ( );
FILL FILL_2_AND2X2_35 ( );
FILL FILL_3_AND2X2_35 ( );
FILL FILL_4_AND2X2_35 ( );
FILL FILL_5_AND2X2_35 ( );
FILL FILL_6_AND2X2_35 ( );
FILL FILL_7_AND2X2_35 ( );
FILL FILL_8_AND2X2_35 ( );
FILL FILL_0_NAND2X1_71 ( );
FILL FILL_1_NAND2X1_71 ( );
FILL FILL_2_NAND2X1_71 ( );
FILL FILL_3_NAND2X1_71 ( );
FILL FILL_4_NAND2X1_71 ( );
FILL FILL_5_NAND2X1_71 ( );
FILL FILL_6_NAND2X1_71 ( );
FILL FILL_0_NAND2X1_81 ( );
FILL FILL_1_NAND2X1_81 ( );
FILL FILL_2_NAND2X1_81 ( );
FILL FILL_3_NAND2X1_81 ( );
FILL FILL_4_NAND2X1_81 ( );
FILL FILL_5_NAND2X1_81 ( );
FILL FILL_6_NAND2X1_81 ( );
FILL FILL_0_NAND3X1_166 ( );
FILL FILL_1_NAND3X1_166 ( );
FILL FILL_2_NAND3X1_166 ( );
FILL FILL_3_NAND3X1_166 ( );
FILL FILL_4_NAND3X1_166 ( );
FILL FILL_5_NAND3X1_166 ( );
FILL FILL_6_NAND3X1_166 ( );
FILL FILL_7_NAND3X1_166 ( );
FILL FILL_8_NAND3X1_166 ( );
FILL FILL_0_OAI21X1_41 ( );
FILL FILL_1_OAI21X1_41 ( );
FILL FILL_2_OAI21X1_41 ( );
FILL FILL_3_OAI21X1_41 ( );
FILL FILL_4_OAI21X1_41 ( );
FILL FILL_5_OAI21X1_41 ( );
FILL FILL_6_OAI21X1_41 ( );
FILL FILL_7_OAI21X1_41 ( );
FILL FILL_8_OAI21X1_41 ( );
FILL FILL_0_AOI21X1_13 ( );
FILL FILL_1_AOI21X1_13 ( );
FILL FILL_2_AOI21X1_13 ( );
FILL FILL_3_AOI21X1_13 ( );
FILL FILL_4_AOI21X1_13 ( );
FILL FILL_5_AOI21X1_13 ( );
FILL FILL_6_AOI21X1_13 ( );
FILL FILL_7_AOI21X1_13 ( );
FILL FILL_8_AOI21X1_13 ( );
FILL FILL_0_OAI21X1_22 ( );
FILL FILL_1_OAI21X1_22 ( );
FILL FILL_2_OAI21X1_22 ( );
FILL FILL_3_OAI21X1_22 ( );
FILL FILL_4_OAI21X1_22 ( );
FILL FILL_5_OAI21X1_22 ( );
FILL FILL_6_OAI21X1_22 ( );
FILL FILL_7_OAI21X1_22 ( );
FILL FILL_8_OAI21X1_22 ( );
FILL FILL_0_AOI21X1_42 ( );
FILL FILL_1_AOI21X1_42 ( );
FILL FILL_2_AOI21X1_42 ( );
FILL FILL_3_AOI21X1_42 ( );
FILL FILL_4_AOI21X1_42 ( );
FILL FILL_5_AOI21X1_42 ( );
FILL FILL_6_AOI21X1_42 ( );
FILL FILL_7_AOI21X1_42 ( );
FILL FILL_8_AOI21X1_42 ( );
FILL FILL_0_NAND2X1_60 ( );
FILL FILL_1_NAND2X1_60 ( );
FILL FILL_2_NAND2X1_60 ( );
FILL FILL_3_NAND2X1_60 ( );
FILL FILL_4_NAND2X1_60 ( );
FILL FILL_5_NAND2X1_60 ( );
FILL FILL_6_NAND2X1_60 ( );
FILL FILL_0_NAND2X1_130 ( );
FILL FILL_1_NAND2X1_130 ( );
FILL FILL_2_NAND2X1_130 ( );
FILL FILL_3_NAND2X1_130 ( );
FILL FILL_4_NAND2X1_130 ( );
FILL FILL_5_NAND2X1_130 ( );
FILL FILL_6_NAND2X1_130 ( );
FILL FILL_0_NAND2X1_135 ( );
FILL FILL_1_NAND2X1_135 ( );
FILL FILL_2_NAND2X1_135 ( );
FILL FILL_3_NAND2X1_135 ( );
FILL FILL_4_NAND2X1_135 ( );
FILL FILL_5_NAND2X1_135 ( );
FILL FILL_6_NAND2X1_135 ( );
FILL FILL_0_OAI21X1_57 ( );
FILL FILL_1_OAI21X1_57 ( );
FILL FILL_2_OAI21X1_57 ( );
FILL FILL_3_OAI21X1_57 ( );
FILL FILL_4_OAI21X1_57 ( );
FILL FILL_5_OAI21X1_57 ( );
FILL FILL_6_OAI21X1_57 ( );
FILL FILL_7_OAI21X1_57 ( );
FILL FILL_8_OAI21X1_57 ( );
FILL FILL_9_OAI21X1_57 ( );
FILL FILL_0_NOR2X1_60 ( );
FILL FILL_1_NOR2X1_60 ( );
FILL FILL_2_NOR2X1_60 ( );
FILL FILL_3_NOR2X1_60 ( );
FILL FILL_4_NOR2X1_60 ( );
FILL FILL_5_NOR2X1_60 ( );
FILL FILL_6_NOR2X1_60 ( );
FILL FILL_0_NAND3X1_130 ( );
FILL FILL_1_NAND3X1_130 ( );
FILL FILL_2_NAND3X1_130 ( );
FILL FILL_3_NAND3X1_130 ( );
FILL FILL_4_NAND3X1_130 ( );
FILL FILL_5_NAND3X1_130 ( );
FILL FILL_6_NAND3X1_130 ( );
FILL FILL_7_NAND3X1_130 ( );
FILL FILL_8_NAND3X1_130 ( );
FILL FILL_9_NAND3X1_130 ( );
FILL FILL_0_AOI21X1_1 ( );
FILL FILL_1_AOI21X1_1 ( );
FILL FILL_2_AOI21X1_1 ( );
FILL FILL_3_AOI21X1_1 ( );
FILL FILL_4_AOI21X1_1 ( );
FILL FILL_5_AOI21X1_1 ( );
FILL FILL_6_AOI21X1_1 ( );
FILL FILL_7_AOI21X1_1 ( );
FILL FILL_8_AOI21X1_1 ( );
FILL FILL_9_AOI21X1_1 ( );
FILL FILL_0_DFFSR_34 ( );
FILL FILL_1_DFFSR_34 ( );
FILL FILL_2_DFFSR_34 ( );
FILL FILL_3_DFFSR_34 ( );
FILL FILL_4_DFFSR_34 ( );
FILL FILL_5_DFFSR_34 ( );
FILL FILL_6_DFFSR_34 ( );
FILL FILL_7_DFFSR_34 ( );
FILL FILL_8_DFFSR_34 ( );
FILL FILL_9_DFFSR_34 ( );
FILL FILL_10_DFFSR_34 ( );
FILL FILL_11_DFFSR_34 ( );
FILL FILL_12_DFFSR_34 ( );
FILL FILL_13_DFFSR_34 ( );
FILL FILL_14_DFFSR_34 ( );
FILL FILL_15_DFFSR_34 ( );
FILL FILL_16_DFFSR_34 ( );
FILL FILL_17_DFFSR_34 ( );
FILL FILL_18_DFFSR_34 ( );
FILL FILL_19_DFFSR_34 ( );
FILL FILL_20_DFFSR_34 ( );
FILL FILL_21_DFFSR_34 ( );
FILL FILL_22_DFFSR_34 ( );
FILL FILL_23_DFFSR_34 ( );
FILL FILL_24_DFFSR_34 ( );
FILL FILL_25_DFFSR_34 ( );
FILL FILL_26_DFFSR_34 ( );
FILL FILL_27_DFFSR_34 ( );
FILL FILL_28_DFFSR_34 ( );
FILL FILL_29_DFFSR_34 ( );
FILL FILL_30_DFFSR_34 ( );
FILL FILL_31_DFFSR_34 ( );
FILL FILL_32_DFFSR_34 ( );
FILL FILL_33_DFFSR_34 ( );
FILL FILL_34_DFFSR_34 ( );
FILL FILL_35_DFFSR_34 ( );
FILL FILL_36_DFFSR_34 ( );
FILL FILL_37_DFFSR_34 ( );
FILL FILL_38_DFFSR_34 ( );
FILL FILL_39_DFFSR_34 ( );
FILL FILL_40_DFFSR_34 ( );
FILL FILL_41_DFFSR_34 ( );
FILL FILL_42_DFFSR_34 ( );
FILL FILL_43_DFFSR_34 ( );
FILL FILL_44_DFFSR_34 ( );
FILL FILL_45_DFFSR_34 ( );
FILL FILL_46_DFFSR_34 ( );
FILL FILL_47_DFFSR_34 ( );
FILL FILL_48_DFFSR_34 ( );
FILL FILL_49_DFFSR_34 ( );
FILL FILL_50_DFFSR_34 ( );
FILL FILL_0_DFFSR_67 ( );
FILL FILL_1_DFFSR_67 ( );
FILL FILL_2_DFFSR_67 ( );
FILL FILL_3_DFFSR_67 ( );
FILL FILL_4_DFFSR_67 ( );
FILL FILL_5_DFFSR_67 ( );
FILL FILL_6_DFFSR_67 ( );
FILL FILL_7_DFFSR_67 ( );
FILL FILL_8_DFFSR_67 ( );
FILL FILL_9_DFFSR_67 ( );
FILL FILL_10_DFFSR_67 ( );
FILL FILL_11_DFFSR_67 ( );
FILL FILL_12_DFFSR_67 ( );
FILL FILL_13_DFFSR_67 ( );
FILL FILL_14_DFFSR_67 ( );
FILL FILL_15_DFFSR_67 ( );
FILL FILL_16_DFFSR_67 ( );
FILL FILL_17_DFFSR_67 ( );
FILL FILL_18_DFFSR_67 ( );
FILL FILL_19_DFFSR_67 ( );
FILL FILL_20_DFFSR_67 ( );
FILL FILL_21_DFFSR_67 ( );
FILL FILL_22_DFFSR_67 ( );
FILL FILL_23_DFFSR_67 ( );
FILL FILL_24_DFFSR_67 ( );
FILL FILL_25_DFFSR_67 ( );
FILL FILL_26_DFFSR_67 ( );
FILL FILL_27_DFFSR_67 ( );
FILL FILL_28_DFFSR_67 ( );
FILL FILL_29_DFFSR_67 ( );
FILL FILL_30_DFFSR_67 ( );
FILL FILL_31_DFFSR_67 ( );
FILL FILL_32_DFFSR_67 ( );
FILL FILL_33_DFFSR_67 ( );
FILL FILL_34_DFFSR_67 ( );
FILL FILL_35_DFFSR_67 ( );
FILL FILL_36_DFFSR_67 ( );
FILL FILL_37_DFFSR_67 ( );
FILL FILL_38_DFFSR_67 ( );
FILL FILL_39_DFFSR_67 ( );
FILL FILL_40_DFFSR_67 ( );
FILL FILL_41_DFFSR_67 ( );
FILL FILL_42_DFFSR_67 ( );
FILL FILL_43_DFFSR_67 ( );
FILL FILL_44_DFFSR_67 ( );
FILL FILL_45_DFFSR_67 ( );
FILL FILL_46_DFFSR_67 ( );
FILL FILL_47_DFFSR_67 ( );
FILL FILL_48_DFFSR_67 ( );
FILL FILL_49_DFFSR_67 ( );
FILL FILL_50_DFFSR_67 ( );
FILL FILL_0_INVX1_181 ( );
FILL FILL_1_INVX1_181 ( );
FILL FILL_2_INVX1_181 ( );
FILL FILL_3_INVX1_181 ( );
FILL FILL_4_INVX1_181 ( );
FILL FILL_0_DFFSR_180 ( );
FILL FILL_1_DFFSR_180 ( );
FILL FILL_2_DFFSR_180 ( );
FILL FILL_3_DFFSR_180 ( );
FILL FILL_4_DFFSR_180 ( );
FILL FILL_5_DFFSR_180 ( );
FILL FILL_6_DFFSR_180 ( );
FILL FILL_7_DFFSR_180 ( );
FILL FILL_8_DFFSR_180 ( );
FILL FILL_9_DFFSR_180 ( );
FILL FILL_10_DFFSR_180 ( );
FILL FILL_11_DFFSR_180 ( );
FILL FILL_12_DFFSR_180 ( );
FILL FILL_13_DFFSR_180 ( );
FILL FILL_14_DFFSR_180 ( );
FILL FILL_15_DFFSR_180 ( );
FILL FILL_16_DFFSR_180 ( );
FILL FILL_17_DFFSR_180 ( );
FILL FILL_18_DFFSR_180 ( );
FILL FILL_19_DFFSR_180 ( );
FILL FILL_20_DFFSR_180 ( );
FILL FILL_21_DFFSR_180 ( );
FILL FILL_22_DFFSR_180 ( );
FILL FILL_23_DFFSR_180 ( );
FILL FILL_24_DFFSR_180 ( );
FILL FILL_25_DFFSR_180 ( );
FILL FILL_26_DFFSR_180 ( );
FILL FILL_27_DFFSR_180 ( );
FILL FILL_28_DFFSR_180 ( );
FILL FILL_29_DFFSR_180 ( );
FILL FILL_30_DFFSR_180 ( );
FILL FILL_31_DFFSR_180 ( );
FILL FILL_32_DFFSR_180 ( );
FILL FILL_33_DFFSR_180 ( );
FILL FILL_34_DFFSR_180 ( );
FILL FILL_35_DFFSR_180 ( );
FILL FILL_36_DFFSR_180 ( );
FILL FILL_37_DFFSR_180 ( );
FILL FILL_38_DFFSR_180 ( );
FILL FILL_39_DFFSR_180 ( );
FILL FILL_40_DFFSR_180 ( );
FILL FILL_41_DFFSR_180 ( );
FILL FILL_42_DFFSR_180 ( );
FILL FILL_43_DFFSR_180 ( );
FILL FILL_44_DFFSR_180 ( );
FILL FILL_45_DFFSR_180 ( );
FILL FILL_46_DFFSR_180 ( );
FILL FILL_47_DFFSR_180 ( );
FILL FILL_48_DFFSR_180 ( );
FILL FILL_49_DFFSR_180 ( );
FILL FILL_50_DFFSR_180 ( );
FILL FILL_0_NOR2X1_43 ( );
FILL FILL_1_NOR2X1_43 ( );
FILL FILL_2_NOR2X1_43 ( );
FILL FILL_3_NOR2X1_43 ( );
FILL FILL_4_NOR2X1_43 ( );
FILL FILL_5_NOR2X1_43 ( );
FILL FILL_6_NOR2X1_43 ( );
FILL FILL_0_NOR2X1_51 ( );
FILL FILL_1_NOR2X1_51 ( );
FILL FILL_2_NOR2X1_51 ( );
FILL FILL_3_NOR2X1_51 ( );
FILL FILL_4_NOR2X1_51 ( );
FILL FILL_5_NOR2X1_51 ( );
FILL FILL_6_NOR2X1_51 ( );
FILL FILL_0_DFFSR_139 ( );
FILL FILL_1_DFFSR_139 ( );
FILL FILL_2_DFFSR_139 ( );
FILL FILL_3_DFFSR_139 ( );
FILL FILL_4_DFFSR_139 ( );
FILL FILL_5_DFFSR_139 ( );
FILL FILL_6_DFFSR_139 ( );
FILL FILL_7_DFFSR_139 ( );
FILL FILL_8_DFFSR_139 ( );
FILL FILL_9_DFFSR_139 ( );
FILL FILL_10_DFFSR_139 ( );
FILL FILL_11_DFFSR_139 ( );
FILL FILL_12_DFFSR_139 ( );
FILL FILL_13_DFFSR_139 ( );
FILL FILL_14_DFFSR_139 ( );
FILL FILL_15_DFFSR_139 ( );
FILL FILL_16_DFFSR_139 ( );
FILL FILL_17_DFFSR_139 ( );
FILL FILL_18_DFFSR_139 ( );
FILL FILL_19_DFFSR_139 ( );
FILL FILL_20_DFFSR_139 ( );
FILL FILL_21_DFFSR_139 ( );
FILL FILL_22_DFFSR_139 ( );
FILL FILL_23_DFFSR_139 ( );
FILL FILL_24_DFFSR_139 ( );
FILL FILL_25_DFFSR_139 ( );
FILL FILL_26_DFFSR_139 ( );
FILL FILL_27_DFFSR_139 ( );
FILL FILL_28_DFFSR_139 ( );
FILL FILL_29_DFFSR_139 ( );
FILL FILL_30_DFFSR_139 ( );
FILL FILL_31_DFFSR_139 ( );
FILL FILL_32_DFFSR_139 ( );
FILL FILL_33_DFFSR_139 ( );
FILL FILL_34_DFFSR_139 ( );
FILL FILL_35_DFFSR_139 ( );
FILL FILL_36_DFFSR_139 ( );
FILL FILL_37_DFFSR_139 ( );
FILL FILL_38_DFFSR_139 ( );
FILL FILL_39_DFFSR_139 ( );
FILL FILL_40_DFFSR_139 ( );
FILL FILL_41_DFFSR_139 ( );
FILL FILL_42_DFFSR_139 ( );
FILL FILL_43_DFFSR_139 ( );
FILL FILL_44_DFFSR_139 ( );
FILL FILL_45_DFFSR_139 ( );
FILL FILL_46_DFFSR_139 ( );
FILL FILL_47_DFFSR_139 ( );
FILL FILL_48_DFFSR_139 ( );
FILL FILL_49_DFFSR_139 ( );
FILL FILL_50_DFFSR_139 ( );
FILL FILL_0_AND2X2_21 ( );
FILL FILL_1_AND2X2_21 ( );
FILL FILL_2_AND2X2_21 ( );
FILL FILL_3_AND2X2_21 ( );
FILL FILL_4_AND2X2_21 ( );
FILL FILL_5_AND2X2_21 ( );
FILL FILL_6_AND2X2_21 ( );
FILL FILL_7_AND2X2_21 ( );
FILL FILL_8_AND2X2_21 ( );
FILL FILL_0_NAND3X1_84 ( );
FILL FILL_1_NAND3X1_84 ( );
FILL FILL_2_NAND3X1_84 ( );
FILL FILL_3_NAND3X1_84 ( );
FILL FILL_4_NAND3X1_84 ( );
FILL FILL_5_NAND3X1_84 ( );
FILL FILL_6_NAND3X1_84 ( );
FILL FILL_7_NAND3X1_84 ( );
FILL FILL_8_NAND3X1_84 ( );
FILL FILL_9_NAND3X1_84 ( );
FILL FILL_0_NOR2X1_32 ( );
FILL FILL_1_NOR2X1_32 ( );
FILL FILL_2_NOR2X1_32 ( );
FILL FILL_3_NOR2X1_32 ( );
FILL FILL_4_NOR2X1_32 ( );
FILL FILL_5_NOR2X1_32 ( );
FILL FILL_6_NOR2X1_32 ( );
FILL FILL_0_NAND2X1_42 ( );
FILL FILL_1_NAND2X1_42 ( );
FILL FILL_2_NAND2X1_42 ( );
FILL FILL_3_NAND2X1_42 ( );
FILL FILL_4_NAND2X1_42 ( );
FILL FILL_5_NAND2X1_42 ( );
FILL FILL_6_NAND2X1_42 ( );
FILL FILL_0_INVX1_107 ( );
FILL FILL_1_INVX1_107 ( );
FILL FILL_2_INVX1_107 ( );
FILL FILL_3_INVX1_107 ( );
FILL FILL_4_INVX1_107 ( );
FILL FILL_0_CLKBUF1_14 ( );
FILL FILL_1_CLKBUF1_14 ( );
FILL FILL_2_CLKBUF1_14 ( );
FILL FILL_3_CLKBUF1_14 ( );
FILL FILL_4_CLKBUF1_14 ( );
FILL FILL_5_CLKBUF1_14 ( );
FILL FILL_6_CLKBUF1_14 ( );
FILL FILL_7_CLKBUF1_14 ( );
FILL FILL_8_CLKBUF1_14 ( );
FILL FILL_9_CLKBUF1_14 ( );
FILL FILL_10_CLKBUF1_14 ( );
FILL FILL_11_CLKBUF1_14 ( );
FILL FILL_12_CLKBUF1_14 ( );
FILL FILL_13_CLKBUF1_14 ( );
FILL FILL_14_CLKBUF1_14 ( );
FILL FILL_15_CLKBUF1_14 ( );
FILL FILL_16_CLKBUF1_14 ( );
FILL FILL_17_CLKBUF1_14 ( );
FILL FILL_18_CLKBUF1_14 ( );
FILL FILL_19_CLKBUF1_14 ( );
FILL FILL_20_CLKBUF1_14 ( );
FILL FILL_0_DFFSR_245 ( );
FILL FILL_1_DFFSR_245 ( );
FILL FILL_2_DFFSR_245 ( );
FILL FILL_3_DFFSR_245 ( );
FILL FILL_4_DFFSR_245 ( );
FILL FILL_5_DFFSR_245 ( );
FILL FILL_6_DFFSR_245 ( );
FILL FILL_7_DFFSR_245 ( );
FILL FILL_8_DFFSR_245 ( );
FILL FILL_9_DFFSR_245 ( );
FILL FILL_10_DFFSR_245 ( );
FILL FILL_11_DFFSR_245 ( );
FILL FILL_12_DFFSR_245 ( );
FILL FILL_13_DFFSR_245 ( );
FILL FILL_14_DFFSR_245 ( );
FILL FILL_15_DFFSR_245 ( );
FILL FILL_16_DFFSR_245 ( );
FILL FILL_17_DFFSR_245 ( );
FILL FILL_18_DFFSR_245 ( );
FILL FILL_19_DFFSR_245 ( );
FILL FILL_20_DFFSR_245 ( );
FILL FILL_21_DFFSR_245 ( );
FILL FILL_22_DFFSR_245 ( );
FILL FILL_23_DFFSR_245 ( );
FILL FILL_24_DFFSR_245 ( );
FILL FILL_25_DFFSR_245 ( );
FILL FILL_26_DFFSR_245 ( );
FILL FILL_27_DFFSR_245 ( );
FILL FILL_28_DFFSR_245 ( );
FILL FILL_29_DFFSR_245 ( );
FILL FILL_30_DFFSR_245 ( );
FILL FILL_31_DFFSR_245 ( );
FILL FILL_32_DFFSR_245 ( );
FILL FILL_33_DFFSR_245 ( );
FILL FILL_34_DFFSR_245 ( );
FILL FILL_35_DFFSR_245 ( );
FILL FILL_36_DFFSR_245 ( );
FILL FILL_37_DFFSR_245 ( );
FILL FILL_38_DFFSR_245 ( );
FILL FILL_39_DFFSR_245 ( );
FILL FILL_40_DFFSR_245 ( );
FILL FILL_41_DFFSR_245 ( );
FILL FILL_42_DFFSR_245 ( );
FILL FILL_43_DFFSR_245 ( );
FILL FILL_44_DFFSR_245 ( );
FILL FILL_45_DFFSR_245 ( );
FILL FILL_46_DFFSR_245 ( );
FILL FILL_47_DFFSR_245 ( );
FILL FILL_48_DFFSR_245 ( );
FILL FILL_49_DFFSR_245 ( );
FILL FILL_50_DFFSR_245 ( );
FILL FILL_51_DFFSR_245 ( );
FILL FILL_0_NAND3X1_182 ( );
FILL FILL_1_NAND3X1_182 ( );
FILL FILL_2_NAND3X1_182 ( );
FILL FILL_3_NAND3X1_182 ( );
FILL FILL_4_NAND3X1_182 ( );
FILL FILL_5_NAND3X1_182 ( );
FILL FILL_6_NAND3X1_182 ( );
FILL FILL_7_NAND3X1_182 ( );
FILL FILL_8_NAND3X1_182 ( );
FILL FILL_9_NAND3X1_182 ( );
FILL FILL_0_NAND2X1_88 ( );
FILL FILL_1_NAND2X1_88 ( );
FILL FILL_2_NAND2X1_88 ( );
FILL FILL_3_NAND2X1_88 ( );
FILL FILL_4_NAND2X1_88 ( );
FILL FILL_5_NAND2X1_88 ( );
FILL FILL_6_NAND2X1_88 ( );
FILL FILL_0_OAI21X1_49 ( );
FILL FILL_1_OAI21X1_49 ( );
FILL FILL_2_OAI21X1_49 ( );
FILL FILL_3_OAI21X1_49 ( );
FILL FILL_4_OAI21X1_49 ( );
FILL FILL_5_OAI21X1_49 ( );
FILL FILL_6_OAI21X1_49 ( );
FILL FILL_7_OAI21X1_49 ( );
FILL FILL_8_OAI21X1_49 ( );
FILL FILL_0_OAI21X1_47 ( );
FILL FILL_1_OAI21X1_47 ( );
FILL FILL_2_OAI21X1_47 ( );
FILL FILL_3_OAI21X1_47 ( );
FILL FILL_4_OAI21X1_47 ( );
FILL FILL_5_OAI21X1_47 ( );
FILL FILL_6_OAI21X1_47 ( );
FILL FILL_7_OAI21X1_47 ( );
FILL FILL_8_OAI21X1_47 ( );
FILL FILL_0_OAI21X1_46 ( );
FILL FILL_1_OAI21X1_46 ( );
FILL FILL_2_OAI21X1_46 ( );
FILL FILL_3_OAI21X1_46 ( );
FILL FILL_4_OAI21X1_46 ( );
FILL FILL_5_OAI21X1_46 ( );
FILL FILL_6_OAI21X1_46 ( );
FILL FILL_7_OAI21X1_46 ( );
FILL FILL_8_OAI21X1_46 ( );
FILL FILL_0_OAI21X1_39 ( );
FILL FILL_1_OAI21X1_39 ( );
FILL FILL_2_OAI21X1_39 ( );
FILL FILL_3_OAI21X1_39 ( );
FILL FILL_4_OAI21X1_39 ( );
FILL FILL_5_OAI21X1_39 ( );
FILL FILL_6_OAI21X1_39 ( );
FILL FILL_7_OAI21X1_39 ( );
FILL FILL_8_OAI21X1_39 ( );
FILL FILL_0_NAND3X1_164 ( );
FILL FILL_1_NAND3X1_164 ( );
FILL FILL_2_NAND3X1_164 ( );
FILL FILL_3_NAND3X1_164 ( );
FILL FILL_4_NAND3X1_164 ( );
FILL FILL_5_NAND3X1_164 ( );
FILL FILL_6_NAND3X1_164 ( );
FILL FILL_7_NAND3X1_164 ( );
FILL FILL_8_NAND3X1_164 ( );
FILL FILL_9_NAND3X1_164 ( );
FILL FILL_0_OAI21X1_40 ( );
FILL FILL_1_OAI21X1_40 ( );
FILL FILL_2_OAI21X1_40 ( );
FILL FILL_3_OAI21X1_40 ( );
FILL FILL_4_OAI21X1_40 ( );
FILL FILL_5_OAI21X1_40 ( );
FILL FILL_6_OAI21X1_40 ( );
FILL FILL_7_OAI21X1_40 ( );
FILL FILL_8_OAI21X1_40 ( );
FILL FILL_0_NAND3X1_152 ( );
FILL FILL_1_NAND3X1_152 ( );
FILL FILL_2_NAND3X1_152 ( );
FILL FILL_3_NAND3X1_152 ( );
FILL FILL_4_NAND3X1_152 ( );
FILL FILL_5_NAND3X1_152 ( );
FILL FILL_6_NAND3X1_152 ( );
FILL FILL_7_NAND3X1_152 ( );
FILL FILL_8_NAND3X1_152 ( );
FILL FILL_0_OAI21X1_24 ( );
FILL FILL_1_OAI21X1_24 ( );
FILL FILL_2_OAI21X1_24 ( );
FILL FILL_3_OAI21X1_24 ( );
FILL FILL_4_OAI21X1_24 ( );
FILL FILL_5_OAI21X1_24 ( );
FILL FILL_6_OAI21X1_24 ( );
FILL FILL_7_OAI21X1_24 ( );
FILL FILL_8_OAI21X1_24 ( );
FILL FILL_9_OAI21X1_24 ( );
FILL FILL_0_OAI21X1_83 ( );
FILL FILL_1_OAI21X1_83 ( );
FILL FILL_2_OAI21X1_83 ( );
FILL FILL_3_OAI21X1_83 ( );
FILL FILL_4_OAI21X1_83 ( );
FILL FILL_5_OAI21X1_83 ( );
FILL FILL_6_OAI21X1_83 ( );
FILL FILL_7_OAI21X1_83 ( );
FILL FILL_8_OAI21X1_83 ( );
FILL FILL_9_OAI21X1_83 ( );
FILL FILL_0_NOR2X1_65 ( );
FILL FILL_1_NOR2X1_65 ( );
FILL FILL_2_NOR2X1_65 ( );
FILL FILL_3_NOR2X1_65 ( );
FILL FILL_4_NOR2X1_65 ( );
FILL FILL_5_NOR2X1_65 ( );
FILL FILL_6_NOR2X1_65 ( );
FILL FILL_0_OAI21X1_99 ( );
FILL FILL_1_OAI21X1_99 ( );
FILL FILL_2_OAI21X1_99 ( );
FILL FILL_3_OAI21X1_99 ( );
FILL FILL_4_OAI21X1_99 ( );
FILL FILL_5_OAI21X1_99 ( );
FILL FILL_6_OAI21X1_99 ( );
FILL FILL_7_OAI21X1_99 ( );
FILL FILL_8_OAI21X1_99 ( );
FILL FILL_9_OAI21X1_99 ( );
FILL FILL_0_INVX1_123 ( );
FILL FILL_1_INVX1_123 ( );
FILL FILL_2_INVX1_123 ( );
FILL FILL_3_INVX1_123 ( );
FILL FILL_0_DFFPOSX1_19 ( );
FILL FILL_1_DFFPOSX1_19 ( );
FILL FILL_2_DFFPOSX1_19 ( );
FILL FILL_3_DFFPOSX1_19 ( );
FILL FILL_4_DFFPOSX1_19 ( );
FILL FILL_5_DFFPOSX1_19 ( );
FILL FILL_6_DFFPOSX1_19 ( );
FILL FILL_7_DFFPOSX1_19 ( );
FILL FILL_8_DFFPOSX1_19 ( );
FILL FILL_9_DFFPOSX1_19 ( );
FILL FILL_10_DFFPOSX1_19 ( );
FILL FILL_11_DFFPOSX1_19 ( );
FILL FILL_12_DFFPOSX1_19 ( );
FILL FILL_13_DFFPOSX1_19 ( );
FILL FILL_14_DFFPOSX1_19 ( );
FILL FILL_15_DFFPOSX1_19 ( );
FILL FILL_16_DFFPOSX1_19 ( );
FILL FILL_17_DFFPOSX1_19 ( );
FILL FILL_18_DFFPOSX1_19 ( );
FILL FILL_19_DFFPOSX1_19 ( );
FILL FILL_20_DFFPOSX1_19 ( );
FILL FILL_21_DFFPOSX1_19 ( );
FILL FILL_22_DFFPOSX1_19 ( );
FILL FILL_23_DFFPOSX1_19 ( );
FILL FILL_24_DFFPOSX1_19 ( );
FILL FILL_25_DFFPOSX1_19 ( );
FILL FILL_26_DFFPOSX1_19 ( );
FILL FILL_27_DFFPOSX1_19 ( );
FILL FILL_0_NOR2X1_59 ( );
FILL FILL_1_NOR2X1_59 ( );
FILL FILL_2_NOR2X1_59 ( );
FILL FILL_3_NOR2X1_59 ( );
FILL FILL_4_NOR2X1_59 ( );
FILL FILL_5_NOR2X1_59 ( );
FILL FILL_6_NOR2X1_59 ( );
FILL FILL_0_INVX1_198 ( );
FILL FILL_1_INVX1_198 ( );
FILL FILL_2_INVX1_198 ( );
FILL FILL_3_INVX1_198 ( );
FILL FILL_0_INVX1_121 ( );
FILL FILL_1_INVX1_121 ( );
FILL FILL_2_INVX1_121 ( );
FILL FILL_3_INVX1_121 ( );
FILL FILL_4_INVX1_121 ( );
FILL FILL_0_DFFPOSX1_27 ( );
FILL FILL_1_DFFPOSX1_27 ( );
FILL FILL_2_DFFPOSX1_27 ( );
FILL FILL_3_DFFPOSX1_27 ( );
FILL FILL_4_DFFPOSX1_27 ( );
FILL FILL_5_DFFPOSX1_27 ( );
FILL FILL_6_DFFPOSX1_27 ( );
FILL FILL_7_DFFPOSX1_27 ( );
FILL FILL_8_DFFPOSX1_27 ( );
FILL FILL_9_DFFPOSX1_27 ( );
FILL FILL_10_DFFPOSX1_27 ( );
FILL FILL_11_DFFPOSX1_27 ( );
FILL FILL_12_DFFPOSX1_27 ( );
FILL FILL_13_DFFPOSX1_27 ( );
FILL FILL_14_DFFPOSX1_27 ( );
FILL FILL_15_DFFPOSX1_27 ( );
FILL FILL_16_DFFPOSX1_27 ( );
FILL FILL_17_DFFPOSX1_27 ( );
FILL FILL_18_DFFPOSX1_27 ( );
FILL FILL_19_DFFPOSX1_27 ( );
FILL FILL_20_DFFPOSX1_27 ( );
FILL FILL_21_DFFPOSX1_27 ( );
FILL FILL_22_DFFPOSX1_27 ( );
FILL FILL_23_DFFPOSX1_27 ( );
FILL FILL_24_DFFPOSX1_27 ( );
FILL FILL_25_DFFPOSX1_27 ( );
FILL FILL_26_DFFPOSX1_27 ( );
FILL FILL_27_DFFPOSX1_27 ( );
FILL FILL_0_INVX1_124 ( );
FILL FILL_1_INVX1_124 ( );
FILL FILL_2_INVX1_124 ( );
FILL FILL_3_INVX1_124 ( );
FILL FILL_0_AOI21X1_3 ( );
FILL FILL_1_AOI21X1_3 ( );
FILL FILL_2_AOI21X1_3 ( );
FILL FILL_3_AOI21X1_3 ( );
FILL FILL_4_AOI21X1_3 ( );
FILL FILL_5_AOI21X1_3 ( );
FILL FILL_6_AOI21X1_3 ( );
FILL FILL_7_AOI21X1_3 ( );
FILL FILL_8_AOI21X1_3 ( );
FILL FILL_9_AOI21X1_3 ( );
FILL FILL_0_DFFSR_75 ( );
FILL FILL_1_DFFSR_75 ( );
FILL FILL_2_DFFSR_75 ( );
FILL FILL_3_DFFSR_75 ( );
FILL FILL_4_DFFSR_75 ( );
FILL FILL_5_DFFSR_75 ( );
FILL FILL_6_DFFSR_75 ( );
FILL FILL_7_DFFSR_75 ( );
FILL FILL_8_DFFSR_75 ( );
FILL FILL_9_DFFSR_75 ( );
FILL FILL_10_DFFSR_75 ( );
FILL FILL_11_DFFSR_75 ( );
FILL FILL_12_DFFSR_75 ( );
FILL FILL_13_DFFSR_75 ( );
FILL FILL_14_DFFSR_75 ( );
FILL FILL_15_DFFSR_75 ( );
FILL FILL_16_DFFSR_75 ( );
FILL FILL_17_DFFSR_75 ( );
FILL FILL_18_DFFSR_75 ( );
FILL FILL_19_DFFSR_75 ( );
FILL FILL_20_DFFSR_75 ( );
FILL FILL_21_DFFSR_75 ( );
FILL FILL_22_DFFSR_75 ( );
FILL FILL_23_DFFSR_75 ( );
FILL FILL_24_DFFSR_75 ( );
FILL FILL_25_DFFSR_75 ( );
FILL FILL_26_DFFSR_75 ( );
FILL FILL_27_DFFSR_75 ( );
FILL FILL_28_DFFSR_75 ( );
FILL FILL_29_DFFSR_75 ( );
FILL FILL_30_DFFSR_75 ( );
FILL FILL_31_DFFSR_75 ( );
FILL FILL_32_DFFSR_75 ( );
FILL FILL_33_DFFSR_75 ( );
FILL FILL_34_DFFSR_75 ( );
FILL FILL_35_DFFSR_75 ( );
FILL FILL_36_DFFSR_75 ( );
FILL FILL_37_DFFSR_75 ( );
FILL FILL_38_DFFSR_75 ( );
FILL FILL_39_DFFSR_75 ( );
FILL FILL_40_DFFSR_75 ( );
FILL FILL_41_DFFSR_75 ( );
FILL FILL_42_DFFSR_75 ( );
FILL FILL_43_DFFSR_75 ( );
FILL FILL_44_DFFSR_75 ( );
FILL FILL_45_DFFSR_75 ( );
FILL FILL_46_DFFSR_75 ( );
FILL FILL_47_DFFSR_75 ( );
FILL FILL_48_DFFSR_75 ( );
FILL FILL_49_DFFSR_75 ( );
FILL FILL_50_DFFSR_75 ( );
FILL FILL_51_DFFSR_75 ( );
FILL FILL_0_OAI22X1_35 ( );
FILL FILL_1_OAI22X1_35 ( );
FILL FILL_2_OAI22X1_35 ( );
FILL FILL_3_OAI22X1_35 ( );
FILL FILL_4_OAI22X1_35 ( );
FILL FILL_5_OAI22X1_35 ( );
FILL FILL_6_OAI22X1_35 ( );
FILL FILL_7_OAI22X1_35 ( );
FILL FILL_8_OAI22X1_35 ( );
FILL FILL_9_OAI22X1_35 ( );
FILL FILL_10_OAI22X1_35 ( );
FILL FILL_11_OAI22X1_35 ( );
FILL FILL_0_OAI22X1_34 ( );
FILL FILL_1_OAI22X1_34 ( );
FILL FILL_2_OAI22X1_34 ( );
FILL FILL_3_OAI22X1_34 ( );
FILL FILL_4_OAI22X1_34 ( );
FILL FILL_5_OAI22X1_34 ( );
FILL FILL_6_OAI22X1_34 ( );
FILL FILL_7_OAI22X1_34 ( );
FILL FILL_8_OAI22X1_34 ( );
FILL FILL_9_OAI22X1_34 ( );
FILL FILL_10_OAI22X1_34 ( );
FILL FILL_11_OAI22X1_34 ( );
FILL FILL_0_NOR2X1_44 ( );
FILL FILL_1_NOR2X1_44 ( );
FILL FILL_2_NOR2X1_44 ( );
FILL FILL_3_NOR2X1_44 ( );
FILL FILL_4_NOR2X1_44 ( );
FILL FILL_5_NOR2X1_44 ( );
FILL FILL_6_NOR2X1_44 ( );
FILL FILL_0_NAND3X1_92 ( );
FILL FILL_1_NAND3X1_92 ( );
FILL FILL_2_NAND3X1_92 ( );
FILL FILL_3_NAND3X1_92 ( );
FILL FILL_4_NAND3X1_92 ( );
FILL FILL_5_NAND3X1_92 ( );
FILL FILL_6_NAND3X1_92 ( );
FILL FILL_7_NAND3X1_92 ( );
FILL FILL_8_NAND3X1_92 ( );
FILL FILL_0_NOR2X1_46 ( );
FILL FILL_1_NOR2X1_46 ( );
FILL FILL_2_NOR2X1_46 ( );
FILL FILL_3_NOR2X1_46 ( );
FILL FILL_4_NOR2X1_46 ( );
FILL FILL_5_NOR2X1_46 ( );
FILL FILL_6_NOR2X1_46 ( );
FILL FILL_0_NAND3X1_96 ( );
FILL FILL_1_NAND3X1_96 ( );
FILL FILL_2_NAND3X1_96 ( );
FILL FILL_3_NAND3X1_96 ( );
FILL FILL_4_NAND3X1_96 ( );
FILL FILL_5_NAND3X1_96 ( );
FILL FILL_6_NAND3X1_96 ( );
FILL FILL_7_NAND3X1_96 ( );
FILL FILL_8_NAND3X1_96 ( );
FILL FILL_0_NOR2X1_45 ( );
FILL FILL_1_NOR2X1_45 ( );
FILL FILL_2_NOR2X1_45 ( );
FILL FILL_3_NOR2X1_45 ( );
FILL FILL_4_NOR2X1_45 ( );
FILL FILL_5_NOR2X1_45 ( );
FILL FILL_6_NOR2X1_45 ( );
FILL FILL_0_DFFSR_254 ( );
FILL FILL_1_DFFSR_254 ( );
FILL FILL_2_DFFSR_254 ( );
FILL FILL_3_DFFSR_254 ( );
FILL FILL_4_DFFSR_254 ( );
FILL FILL_5_DFFSR_254 ( );
FILL FILL_6_DFFSR_254 ( );
FILL FILL_7_DFFSR_254 ( );
FILL FILL_8_DFFSR_254 ( );
FILL FILL_9_DFFSR_254 ( );
FILL FILL_10_DFFSR_254 ( );
FILL FILL_11_DFFSR_254 ( );
FILL FILL_12_DFFSR_254 ( );
FILL FILL_13_DFFSR_254 ( );
FILL FILL_14_DFFSR_254 ( );
FILL FILL_15_DFFSR_254 ( );
FILL FILL_16_DFFSR_254 ( );
FILL FILL_17_DFFSR_254 ( );
FILL FILL_18_DFFSR_254 ( );
FILL FILL_19_DFFSR_254 ( );
FILL FILL_20_DFFSR_254 ( );
FILL FILL_21_DFFSR_254 ( );
FILL FILL_22_DFFSR_254 ( );
FILL FILL_23_DFFSR_254 ( );
FILL FILL_24_DFFSR_254 ( );
FILL FILL_25_DFFSR_254 ( );
FILL FILL_26_DFFSR_254 ( );
FILL FILL_27_DFFSR_254 ( );
FILL FILL_28_DFFSR_254 ( );
FILL FILL_29_DFFSR_254 ( );
FILL FILL_30_DFFSR_254 ( );
FILL FILL_31_DFFSR_254 ( );
FILL FILL_32_DFFSR_254 ( );
FILL FILL_33_DFFSR_254 ( );
FILL FILL_34_DFFSR_254 ( );
FILL FILL_35_DFFSR_254 ( );
FILL FILL_36_DFFSR_254 ( );
FILL FILL_37_DFFSR_254 ( );
FILL FILL_38_DFFSR_254 ( );
FILL FILL_39_DFFSR_254 ( );
FILL FILL_40_DFFSR_254 ( );
FILL FILL_41_DFFSR_254 ( );
FILL FILL_42_DFFSR_254 ( );
FILL FILL_43_DFFSR_254 ( );
FILL FILL_44_DFFSR_254 ( );
FILL FILL_45_DFFSR_254 ( );
FILL FILL_46_DFFSR_254 ( );
FILL FILL_47_DFFSR_254 ( );
FILL FILL_48_DFFSR_254 ( );
FILL FILL_49_DFFSR_254 ( );
FILL FILL_50_DFFSR_254 ( );
FILL FILL_51_DFFSR_254 ( );
FILL FILL_0_DFFSR_215 ( );
FILL FILL_1_DFFSR_215 ( );
FILL FILL_2_DFFSR_215 ( );
FILL FILL_3_DFFSR_215 ( );
FILL FILL_4_DFFSR_215 ( );
FILL FILL_5_DFFSR_215 ( );
FILL FILL_6_DFFSR_215 ( );
FILL FILL_7_DFFSR_215 ( );
FILL FILL_8_DFFSR_215 ( );
FILL FILL_9_DFFSR_215 ( );
FILL FILL_10_DFFSR_215 ( );
FILL FILL_11_DFFSR_215 ( );
FILL FILL_12_DFFSR_215 ( );
FILL FILL_13_DFFSR_215 ( );
FILL FILL_14_DFFSR_215 ( );
FILL FILL_15_DFFSR_215 ( );
FILL FILL_16_DFFSR_215 ( );
FILL FILL_17_DFFSR_215 ( );
FILL FILL_18_DFFSR_215 ( );
FILL FILL_19_DFFSR_215 ( );
FILL FILL_20_DFFSR_215 ( );
FILL FILL_21_DFFSR_215 ( );
FILL FILL_22_DFFSR_215 ( );
FILL FILL_23_DFFSR_215 ( );
FILL FILL_24_DFFSR_215 ( );
FILL FILL_25_DFFSR_215 ( );
FILL FILL_26_DFFSR_215 ( );
FILL FILL_27_DFFSR_215 ( );
FILL FILL_28_DFFSR_215 ( );
FILL FILL_29_DFFSR_215 ( );
FILL FILL_30_DFFSR_215 ( );
FILL FILL_31_DFFSR_215 ( );
FILL FILL_32_DFFSR_215 ( );
FILL FILL_33_DFFSR_215 ( );
FILL FILL_34_DFFSR_215 ( );
FILL FILL_35_DFFSR_215 ( );
FILL FILL_36_DFFSR_215 ( );
FILL FILL_37_DFFSR_215 ( );
FILL FILL_38_DFFSR_215 ( );
FILL FILL_39_DFFSR_215 ( );
FILL FILL_40_DFFSR_215 ( );
FILL FILL_41_DFFSR_215 ( );
FILL FILL_42_DFFSR_215 ( );
FILL FILL_43_DFFSR_215 ( );
FILL FILL_44_DFFSR_215 ( );
FILL FILL_45_DFFSR_215 ( );
FILL FILL_46_DFFSR_215 ( );
FILL FILL_47_DFFSR_215 ( );
FILL FILL_48_DFFSR_215 ( );
FILL FILL_49_DFFSR_215 ( );
FILL FILL_50_DFFSR_215 ( );
FILL FILL_0_DFFSR_253 ( );
FILL FILL_1_DFFSR_253 ( );
FILL FILL_2_DFFSR_253 ( );
FILL FILL_3_DFFSR_253 ( );
FILL FILL_4_DFFSR_253 ( );
FILL FILL_5_DFFSR_253 ( );
FILL FILL_6_DFFSR_253 ( );
FILL FILL_7_DFFSR_253 ( );
FILL FILL_8_DFFSR_253 ( );
FILL FILL_9_DFFSR_253 ( );
FILL FILL_10_DFFSR_253 ( );
FILL FILL_11_DFFSR_253 ( );
FILL FILL_12_DFFSR_253 ( );
FILL FILL_13_DFFSR_253 ( );
FILL FILL_14_DFFSR_253 ( );
FILL FILL_15_DFFSR_253 ( );
FILL FILL_16_DFFSR_253 ( );
FILL FILL_17_DFFSR_253 ( );
FILL FILL_18_DFFSR_253 ( );
FILL FILL_19_DFFSR_253 ( );
FILL FILL_20_DFFSR_253 ( );
FILL FILL_21_DFFSR_253 ( );
FILL FILL_22_DFFSR_253 ( );
FILL FILL_23_DFFSR_253 ( );
FILL FILL_24_DFFSR_253 ( );
FILL FILL_25_DFFSR_253 ( );
FILL FILL_26_DFFSR_253 ( );
FILL FILL_27_DFFSR_253 ( );
FILL FILL_28_DFFSR_253 ( );
FILL FILL_29_DFFSR_253 ( );
FILL FILL_30_DFFSR_253 ( );
FILL FILL_31_DFFSR_253 ( );
FILL FILL_32_DFFSR_253 ( );
FILL FILL_33_DFFSR_253 ( );
FILL FILL_34_DFFSR_253 ( );
FILL FILL_35_DFFSR_253 ( );
FILL FILL_36_DFFSR_253 ( );
FILL FILL_37_DFFSR_253 ( );
FILL FILL_38_DFFSR_253 ( );
FILL FILL_39_DFFSR_253 ( );
FILL FILL_40_DFFSR_253 ( );
FILL FILL_41_DFFSR_253 ( );
FILL FILL_42_DFFSR_253 ( );
FILL FILL_43_DFFSR_253 ( );
FILL FILL_44_DFFSR_253 ( );
FILL FILL_45_DFFSR_253 ( );
FILL FILL_46_DFFSR_253 ( );
FILL FILL_47_DFFSR_253 ( );
FILL FILL_48_DFFSR_253 ( );
FILL FILL_49_DFFSR_253 ( );
FILL FILL_50_DFFSR_253 ( );
FILL FILL_0_NAND3X1_172 ( );
FILL FILL_1_NAND3X1_172 ( );
FILL FILL_2_NAND3X1_172 ( );
FILL FILL_3_NAND3X1_172 ( );
FILL FILL_4_NAND3X1_172 ( );
FILL FILL_5_NAND3X1_172 ( );
FILL FILL_6_NAND3X1_172 ( );
FILL FILL_7_NAND3X1_172 ( );
FILL FILL_8_NAND3X1_172 ( );
FILL FILL_9_NAND3X1_172 ( );
FILL FILL_0_OAI21X1_61 ( );
FILL FILL_1_OAI21X1_61 ( );
FILL FILL_2_OAI21X1_61 ( );
FILL FILL_3_OAI21X1_61 ( );
FILL FILL_4_OAI21X1_61 ( );
FILL FILL_5_OAI21X1_61 ( );
FILL FILL_6_OAI21X1_61 ( );
FILL FILL_7_OAI21X1_61 ( );
FILL FILL_8_OAI21X1_61 ( );
FILL FILL_0_NAND3X1_207 ( );
FILL FILL_1_NAND3X1_207 ( );
FILL FILL_2_NAND3X1_207 ( );
FILL FILL_3_NAND3X1_207 ( );
FILL FILL_4_NAND3X1_207 ( );
FILL FILL_5_NAND3X1_207 ( );
FILL FILL_6_NAND3X1_207 ( );
FILL FILL_7_NAND3X1_207 ( );
FILL FILL_8_NAND3X1_207 ( );
FILL FILL_0_AOI21X1_20 ( );
FILL FILL_1_AOI21X1_20 ( );
FILL FILL_2_AOI21X1_20 ( );
FILL FILL_3_AOI21X1_20 ( );
FILL FILL_4_AOI21X1_20 ( );
FILL FILL_5_AOI21X1_20 ( );
FILL FILL_6_AOI21X1_20 ( );
FILL FILL_7_AOI21X1_20 ( );
FILL FILL_8_AOI21X1_20 ( );
FILL FILL_9_AOI21X1_20 ( );
FILL FILL_0_NAND3X1_163 ( );
FILL FILL_1_NAND3X1_163 ( );
FILL FILL_2_NAND3X1_163 ( );
FILL FILL_3_NAND3X1_163 ( );
FILL FILL_4_NAND3X1_163 ( );
FILL FILL_5_NAND3X1_163 ( );
FILL FILL_6_NAND3X1_163 ( );
FILL FILL_7_NAND3X1_163 ( );
FILL FILL_8_NAND3X1_163 ( );
FILL FILL_0_NAND3X1_149 ( );
FILL FILL_1_NAND3X1_149 ( );
FILL FILL_2_NAND3X1_149 ( );
FILL FILL_3_NAND3X1_149 ( );
FILL FILL_4_NAND3X1_149 ( );
FILL FILL_5_NAND3X1_149 ( );
FILL FILL_6_NAND3X1_149 ( );
FILL FILL_7_NAND3X1_149 ( );
FILL FILL_8_NAND3X1_149 ( );
FILL FILL_0_AOI21X1_12 ( );
FILL FILL_1_AOI21X1_12 ( );
FILL FILL_2_AOI21X1_12 ( );
FILL FILL_3_AOI21X1_12 ( );
FILL FILL_4_AOI21X1_12 ( );
FILL FILL_5_AOI21X1_12 ( );
FILL FILL_6_AOI21X1_12 ( );
FILL FILL_7_AOI21X1_12 ( );
FILL FILL_8_AOI21X1_12 ( );
FILL FILL_0_NAND3X1_150 ( );
FILL FILL_1_NAND3X1_150 ( );
FILL FILL_2_NAND3X1_150 ( );
FILL FILL_3_NAND3X1_150 ( );
FILL FILL_4_NAND3X1_150 ( );
FILL FILL_5_NAND3X1_150 ( );
FILL FILL_6_NAND3X1_150 ( );
FILL FILL_7_NAND3X1_150 ( );
FILL FILL_8_NAND3X1_150 ( );
FILL FILL_0_NAND3X1_140 ( );
FILL FILL_1_NAND3X1_140 ( );
FILL FILL_2_NAND3X1_140 ( );
FILL FILL_3_NAND3X1_140 ( );
FILL FILL_4_NAND3X1_140 ( );
FILL FILL_5_NAND3X1_140 ( );
FILL FILL_6_NAND3X1_140 ( );
FILL FILL_7_NAND3X1_140 ( );
FILL FILL_8_NAND3X1_140 ( );
FILL FILL_0_AOI21X1_8 ( );
FILL FILL_1_AOI21X1_8 ( );
FILL FILL_2_AOI21X1_8 ( );
FILL FILL_3_AOI21X1_8 ( );
FILL FILL_4_AOI21X1_8 ( );
FILL FILL_5_AOI21X1_8 ( );
FILL FILL_6_AOI21X1_8 ( );
FILL FILL_7_AOI21X1_8 ( );
FILL FILL_8_AOI21X1_8 ( );
FILL FILL_9_AOI21X1_8 ( );
FILL FILL_0_BUFX2_55 ( );
FILL FILL_1_BUFX2_55 ( );
FILL FILL_2_BUFX2_55 ( );
FILL FILL_3_BUFX2_55 ( );
FILL FILL_4_BUFX2_55 ( );
FILL FILL_5_BUFX2_55 ( );
FILL FILL_6_BUFX2_55 ( );
FILL FILL_0_NAND2X1_134 ( );
FILL FILL_1_NAND2X1_134 ( );
FILL FILL_2_NAND2X1_134 ( );
FILL FILL_3_NAND2X1_134 ( );
FILL FILL_4_NAND2X1_134 ( );
FILL FILL_5_NAND2X1_134 ( );
FILL FILL_6_NAND2X1_134 ( );
FILL FILL_0_BUFX2_38 ( );
FILL FILL_1_BUFX2_38 ( );
FILL FILL_2_BUFX2_38 ( );
FILL FILL_3_BUFX2_38 ( );
FILL FILL_4_BUFX2_38 ( );
FILL FILL_5_BUFX2_38 ( );
FILL FILL_6_BUFX2_38 ( );
FILL FILL_0_INVX1_207 ( );
FILL FILL_1_INVX1_207 ( );
FILL FILL_2_INVX1_207 ( );
FILL FILL_3_INVX1_207 ( );
FILL FILL_4_INVX1_207 ( );
FILL FILL_0_INVX1_122 ( );
FILL FILL_1_INVX1_122 ( );
FILL FILL_2_INVX1_122 ( );
FILL FILL_3_INVX1_122 ( );
FILL FILL_4_INVX1_122 ( );
FILL FILL_0_DFFPOSX1_2 ( );
FILL FILL_1_DFFPOSX1_2 ( );
FILL FILL_2_DFFPOSX1_2 ( );
FILL FILL_3_DFFPOSX1_2 ( );
FILL FILL_4_DFFPOSX1_2 ( );
FILL FILL_5_DFFPOSX1_2 ( );
FILL FILL_6_DFFPOSX1_2 ( );
FILL FILL_7_DFFPOSX1_2 ( );
FILL FILL_8_DFFPOSX1_2 ( );
FILL FILL_9_DFFPOSX1_2 ( );
FILL FILL_10_DFFPOSX1_2 ( );
FILL FILL_11_DFFPOSX1_2 ( );
FILL FILL_12_DFFPOSX1_2 ( );
FILL FILL_13_DFFPOSX1_2 ( );
FILL FILL_14_DFFPOSX1_2 ( );
FILL FILL_15_DFFPOSX1_2 ( );
FILL FILL_16_DFFPOSX1_2 ( );
FILL FILL_17_DFFPOSX1_2 ( );
FILL FILL_18_DFFPOSX1_2 ( );
FILL FILL_19_DFFPOSX1_2 ( );
FILL FILL_20_DFFPOSX1_2 ( );
FILL FILL_21_DFFPOSX1_2 ( );
FILL FILL_22_DFFPOSX1_2 ( );
FILL FILL_23_DFFPOSX1_2 ( );
FILL FILL_24_DFFPOSX1_2 ( );
FILL FILL_25_DFFPOSX1_2 ( );
FILL FILL_26_DFFPOSX1_2 ( );
FILL FILL_27_DFFPOSX1_2 ( );
FILL FILL_0_NAND2X1_150 ( );
FILL FILL_1_NAND2X1_150 ( );
FILL FILL_2_NAND2X1_150 ( );
FILL FILL_3_NAND2X1_150 ( );
FILL FILL_4_NAND2X1_150 ( );
FILL FILL_5_NAND2X1_150 ( );
FILL FILL_6_NAND2X1_150 ( );
FILL FILL_0_NAND2X1_57 ( );
FILL FILL_1_NAND2X1_57 ( );
FILL FILL_2_NAND2X1_57 ( );
FILL FILL_3_NAND2X1_57 ( );
FILL FILL_4_NAND2X1_57 ( );
FILL FILL_5_NAND2X1_57 ( );
FILL FILL_6_NAND2X1_57 ( );
FILL FILL_0_DFFSR_11 ( );
FILL FILL_1_DFFSR_11 ( );
FILL FILL_2_DFFSR_11 ( );
FILL FILL_3_DFFSR_11 ( );
FILL FILL_4_DFFSR_11 ( );
FILL FILL_5_DFFSR_11 ( );
FILL FILL_6_DFFSR_11 ( );
FILL FILL_7_DFFSR_11 ( );
FILL FILL_8_DFFSR_11 ( );
FILL FILL_9_DFFSR_11 ( );
FILL FILL_10_DFFSR_11 ( );
FILL FILL_11_DFFSR_11 ( );
FILL FILL_12_DFFSR_11 ( );
FILL FILL_13_DFFSR_11 ( );
FILL FILL_14_DFFSR_11 ( );
FILL FILL_15_DFFSR_11 ( );
FILL FILL_16_DFFSR_11 ( );
FILL FILL_17_DFFSR_11 ( );
FILL FILL_18_DFFSR_11 ( );
FILL FILL_19_DFFSR_11 ( );
FILL FILL_20_DFFSR_11 ( );
FILL FILL_21_DFFSR_11 ( );
FILL FILL_22_DFFSR_11 ( );
FILL FILL_23_DFFSR_11 ( );
FILL FILL_24_DFFSR_11 ( );
FILL FILL_25_DFFSR_11 ( );
FILL FILL_26_DFFSR_11 ( );
FILL FILL_27_DFFSR_11 ( );
FILL FILL_28_DFFSR_11 ( );
FILL FILL_29_DFFSR_11 ( );
FILL FILL_30_DFFSR_11 ( );
FILL FILL_31_DFFSR_11 ( );
FILL FILL_32_DFFSR_11 ( );
FILL FILL_33_DFFSR_11 ( );
FILL FILL_34_DFFSR_11 ( );
FILL FILL_35_DFFSR_11 ( );
FILL FILL_36_DFFSR_11 ( );
FILL FILL_37_DFFSR_11 ( );
FILL FILL_38_DFFSR_11 ( );
FILL FILL_39_DFFSR_11 ( );
FILL FILL_40_DFFSR_11 ( );
FILL FILL_41_DFFSR_11 ( );
FILL FILL_42_DFFSR_11 ( );
FILL FILL_43_DFFSR_11 ( );
FILL FILL_44_DFFSR_11 ( );
FILL FILL_45_DFFSR_11 ( );
FILL FILL_46_DFFSR_11 ( );
FILL FILL_47_DFFSR_11 ( );
FILL FILL_48_DFFSR_11 ( );
FILL FILL_49_DFFSR_11 ( );
FILL FILL_50_DFFSR_11 ( );
FILL FILL_51_DFFSR_11 ( );
FILL FILL_0_DFFSR_1 ( );
FILL FILL_1_DFFSR_1 ( );
FILL FILL_2_DFFSR_1 ( );
FILL FILL_3_DFFSR_1 ( );
FILL FILL_4_DFFSR_1 ( );
FILL FILL_5_DFFSR_1 ( );
FILL FILL_6_DFFSR_1 ( );
FILL FILL_7_DFFSR_1 ( );
FILL FILL_8_DFFSR_1 ( );
FILL FILL_9_DFFSR_1 ( );
FILL FILL_10_DFFSR_1 ( );
FILL FILL_11_DFFSR_1 ( );
FILL FILL_12_DFFSR_1 ( );
FILL FILL_13_DFFSR_1 ( );
FILL FILL_14_DFFSR_1 ( );
FILL FILL_15_DFFSR_1 ( );
FILL FILL_16_DFFSR_1 ( );
FILL FILL_17_DFFSR_1 ( );
FILL FILL_18_DFFSR_1 ( );
FILL FILL_19_DFFSR_1 ( );
FILL FILL_20_DFFSR_1 ( );
FILL FILL_21_DFFSR_1 ( );
FILL FILL_22_DFFSR_1 ( );
FILL FILL_23_DFFSR_1 ( );
FILL FILL_24_DFFSR_1 ( );
FILL FILL_25_DFFSR_1 ( );
FILL FILL_26_DFFSR_1 ( );
FILL FILL_27_DFFSR_1 ( );
FILL FILL_28_DFFSR_1 ( );
FILL FILL_29_DFFSR_1 ( );
FILL FILL_30_DFFSR_1 ( );
FILL FILL_31_DFFSR_1 ( );
FILL FILL_32_DFFSR_1 ( );
FILL FILL_33_DFFSR_1 ( );
FILL FILL_34_DFFSR_1 ( );
FILL FILL_35_DFFSR_1 ( );
FILL FILL_36_DFFSR_1 ( );
FILL FILL_37_DFFSR_1 ( );
FILL FILL_38_DFFSR_1 ( );
FILL FILL_39_DFFSR_1 ( );
FILL FILL_40_DFFSR_1 ( );
FILL FILL_41_DFFSR_1 ( );
FILL FILL_42_DFFSR_1 ( );
FILL FILL_43_DFFSR_1 ( );
FILL FILL_44_DFFSR_1 ( );
FILL FILL_45_DFFSR_1 ( );
FILL FILL_46_DFFSR_1 ( );
FILL FILL_47_DFFSR_1 ( );
FILL FILL_48_DFFSR_1 ( );
FILL FILL_49_DFFSR_1 ( );
FILL FILL_50_DFFSR_1 ( );
FILL FILL_0_NAND3X1_112 ( );
FILL FILL_1_NAND3X1_112 ( );
FILL FILL_2_NAND3X1_112 ( );
FILL FILL_3_NAND3X1_112 ( );
FILL FILL_4_NAND3X1_112 ( );
FILL FILL_5_NAND3X1_112 ( );
FILL FILL_6_NAND3X1_112 ( );
FILL FILL_7_NAND3X1_112 ( );
FILL FILL_8_NAND3X1_112 ( );
FILL FILL_9_NAND3X1_112 ( );
FILL FILL_0_NOR2X1_52 ( );
FILL FILL_1_NOR2X1_52 ( );
FILL FILL_2_NOR2X1_52 ( );
FILL FILL_3_NOR2X1_52 ( );
FILL FILL_4_NOR2X1_52 ( );
FILL FILL_5_NOR2X1_52 ( );
FILL FILL_6_NOR2X1_52 ( );
FILL FILL_0_DFFSR_147 ( );
FILL FILL_1_DFFSR_147 ( );
FILL FILL_2_DFFSR_147 ( );
FILL FILL_3_DFFSR_147 ( );
FILL FILL_4_DFFSR_147 ( );
FILL FILL_5_DFFSR_147 ( );
FILL FILL_6_DFFSR_147 ( );
FILL FILL_7_DFFSR_147 ( );
FILL FILL_8_DFFSR_147 ( );
FILL FILL_9_DFFSR_147 ( );
FILL FILL_10_DFFSR_147 ( );
FILL FILL_11_DFFSR_147 ( );
FILL FILL_12_DFFSR_147 ( );
FILL FILL_13_DFFSR_147 ( );
FILL FILL_14_DFFSR_147 ( );
FILL FILL_15_DFFSR_147 ( );
FILL FILL_16_DFFSR_147 ( );
FILL FILL_17_DFFSR_147 ( );
FILL FILL_18_DFFSR_147 ( );
FILL FILL_19_DFFSR_147 ( );
FILL FILL_20_DFFSR_147 ( );
FILL FILL_21_DFFSR_147 ( );
FILL FILL_22_DFFSR_147 ( );
FILL FILL_23_DFFSR_147 ( );
FILL FILL_24_DFFSR_147 ( );
FILL FILL_25_DFFSR_147 ( );
FILL FILL_26_DFFSR_147 ( );
FILL FILL_27_DFFSR_147 ( );
FILL FILL_28_DFFSR_147 ( );
FILL FILL_29_DFFSR_147 ( );
FILL FILL_30_DFFSR_147 ( );
FILL FILL_31_DFFSR_147 ( );
FILL FILL_32_DFFSR_147 ( );
FILL FILL_33_DFFSR_147 ( );
FILL FILL_34_DFFSR_147 ( );
FILL FILL_35_DFFSR_147 ( );
FILL FILL_36_DFFSR_147 ( );
FILL FILL_37_DFFSR_147 ( );
FILL FILL_38_DFFSR_147 ( );
FILL FILL_39_DFFSR_147 ( );
FILL FILL_40_DFFSR_147 ( );
FILL FILL_41_DFFSR_147 ( );
FILL FILL_42_DFFSR_147 ( );
FILL FILL_43_DFFSR_147 ( );
FILL FILL_44_DFFSR_147 ( );
FILL FILL_45_DFFSR_147 ( );
FILL FILL_46_DFFSR_147 ( );
FILL FILL_47_DFFSR_147 ( );
FILL FILL_48_DFFSR_147 ( );
FILL FILL_49_DFFSR_147 ( );
FILL FILL_50_DFFSR_147 ( );
FILL FILL_0_INVX1_76 ( );
FILL FILL_1_INVX1_76 ( );
FILL FILL_2_INVX1_76 ( );
FILL FILL_3_INVX1_76 ( );
FILL FILL_4_INVX1_76 ( );
FILL FILL_0_BUFX2_69 ( );
FILL FILL_1_BUFX2_69 ( );
FILL FILL_2_BUFX2_69 ( );
FILL FILL_3_BUFX2_69 ( );
FILL FILL_4_BUFX2_69 ( );
FILL FILL_5_BUFX2_69 ( );
FILL FILL_6_BUFX2_69 ( );
FILL FILL_0_NAND3X1_82 ( );
FILL FILL_1_NAND3X1_82 ( );
FILL FILL_2_NAND3X1_82 ( );
FILL FILL_3_NAND3X1_82 ( );
FILL FILL_4_NAND3X1_82 ( );
FILL FILL_5_NAND3X1_82 ( );
FILL FILL_6_NAND3X1_82 ( );
FILL FILL_7_NAND3X1_82 ( );
FILL FILL_8_NAND3X1_82 ( );
FILL FILL_9_NAND3X1_82 ( );
FILL FILL_0_NAND3X1_81 ( );
FILL FILL_1_NAND3X1_81 ( );
FILL FILL_2_NAND3X1_81 ( );
FILL FILL_3_NAND3X1_81 ( );
FILL FILL_4_NAND3X1_81 ( );
FILL FILL_5_NAND3X1_81 ( );
FILL FILL_6_NAND3X1_81 ( );
FILL FILL_7_NAND3X1_81 ( );
FILL FILL_8_NAND3X1_81 ( );
FILL FILL_0_DFFSR_163 ( );
FILL FILL_1_DFFSR_163 ( );
FILL FILL_2_DFFSR_163 ( );
FILL FILL_3_DFFSR_163 ( );
FILL FILL_4_DFFSR_163 ( );
FILL FILL_5_DFFSR_163 ( );
FILL FILL_6_DFFSR_163 ( );
FILL FILL_7_DFFSR_163 ( );
FILL FILL_8_DFFSR_163 ( );
FILL FILL_9_DFFSR_163 ( );
FILL FILL_10_DFFSR_163 ( );
FILL FILL_11_DFFSR_163 ( );
FILL FILL_12_DFFSR_163 ( );
FILL FILL_13_DFFSR_163 ( );
FILL FILL_14_DFFSR_163 ( );
FILL FILL_15_DFFSR_163 ( );
FILL FILL_16_DFFSR_163 ( );
FILL FILL_17_DFFSR_163 ( );
FILL FILL_18_DFFSR_163 ( );
FILL FILL_19_DFFSR_163 ( );
FILL FILL_20_DFFSR_163 ( );
FILL FILL_21_DFFSR_163 ( );
FILL FILL_22_DFFSR_163 ( );
FILL FILL_23_DFFSR_163 ( );
FILL FILL_24_DFFSR_163 ( );
FILL FILL_25_DFFSR_163 ( );
FILL FILL_26_DFFSR_163 ( );
FILL FILL_27_DFFSR_163 ( );
FILL FILL_28_DFFSR_163 ( );
FILL FILL_29_DFFSR_163 ( );
FILL FILL_30_DFFSR_163 ( );
FILL FILL_31_DFFSR_163 ( );
FILL FILL_32_DFFSR_163 ( );
FILL FILL_33_DFFSR_163 ( );
FILL FILL_34_DFFSR_163 ( );
FILL FILL_35_DFFSR_163 ( );
FILL FILL_36_DFFSR_163 ( );
FILL FILL_37_DFFSR_163 ( );
FILL FILL_38_DFFSR_163 ( );
FILL FILL_39_DFFSR_163 ( );
FILL FILL_40_DFFSR_163 ( );
FILL FILL_41_DFFSR_163 ( );
FILL FILL_42_DFFSR_163 ( );
FILL FILL_43_DFFSR_163 ( );
FILL FILL_44_DFFSR_163 ( );
FILL FILL_45_DFFSR_163 ( );
FILL FILL_46_DFFSR_163 ( );
FILL FILL_47_DFFSR_163 ( );
FILL FILL_48_DFFSR_163 ( );
FILL FILL_49_DFFSR_163 ( );
FILL FILL_50_DFFSR_163 ( );
FILL FILL_0_INVX1_73 ( );
FILL FILL_1_INVX1_73 ( );
FILL FILL_2_INVX1_73 ( );
FILL FILL_3_INVX1_73 ( );
FILL FILL_4_INVX1_73 ( );
FILL FILL_0_DFFSR_237 ( );
FILL FILL_1_DFFSR_237 ( );
FILL FILL_2_DFFSR_237 ( );
FILL FILL_3_DFFSR_237 ( );
FILL FILL_4_DFFSR_237 ( );
FILL FILL_5_DFFSR_237 ( );
FILL FILL_6_DFFSR_237 ( );
FILL FILL_7_DFFSR_237 ( );
FILL FILL_8_DFFSR_237 ( );
FILL FILL_9_DFFSR_237 ( );
FILL FILL_10_DFFSR_237 ( );
FILL FILL_11_DFFSR_237 ( );
FILL FILL_12_DFFSR_237 ( );
FILL FILL_13_DFFSR_237 ( );
FILL FILL_14_DFFSR_237 ( );
FILL FILL_15_DFFSR_237 ( );
FILL FILL_16_DFFSR_237 ( );
FILL FILL_17_DFFSR_237 ( );
FILL FILL_18_DFFSR_237 ( );
FILL FILL_19_DFFSR_237 ( );
FILL FILL_20_DFFSR_237 ( );
FILL FILL_21_DFFSR_237 ( );
FILL FILL_22_DFFSR_237 ( );
FILL FILL_23_DFFSR_237 ( );
FILL FILL_24_DFFSR_237 ( );
FILL FILL_25_DFFSR_237 ( );
FILL FILL_26_DFFSR_237 ( );
FILL FILL_27_DFFSR_237 ( );
FILL FILL_28_DFFSR_237 ( );
FILL FILL_29_DFFSR_237 ( );
FILL FILL_30_DFFSR_237 ( );
FILL FILL_31_DFFSR_237 ( );
FILL FILL_32_DFFSR_237 ( );
FILL FILL_33_DFFSR_237 ( );
FILL FILL_34_DFFSR_237 ( );
FILL FILL_35_DFFSR_237 ( );
FILL FILL_36_DFFSR_237 ( );
FILL FILL_37_DFFSR_237 ( );
FILL FILL_38_DFFSR_237 ( );
FILL FILL_39_DFFSR_237 ( );
FILL FILL_40_DFFSR_237 ( );
FILL FILL_41_DFFSR_237 ( );
FILL FILL_42_DFFSR_237 ( );
FILL FILL_43_DFFSR_237 ( );
FILL FILL_44_DFFSR_237 ( );
FILL FILL_45_DFFSR_237 ( );
FILL FILL_46_DFFSR_237 ( );
FILL FILL_47_DFFSR_237 ( );
FILL FILL_48_DFFSR_237 ( );
FILL FILL_49_DFFSR_237 ( );
FILL FILL_50_DFFSR_237 ( );
FILL FILL_0_NAND2X1_82 ( );
FILL FILL_1_NAND2X1_82 ( );
FILL FILL_2_NAND2X1_82 ( );
FILL FILL_3_NAND2X1_82 ( );
FILL FILL_4_NAND2X1_82 ( );
FILL FILL_5_NAND2X1_82 ( );
FILL FILL_6_NAND2X1_82 ( );
FILL FILL_0_NAND3X1_211 ( );
FILL FILL_1_NAND3X1_211 ( );
FILL FILL_2_NAND3X1_211 ( );
FILL FILL_3_NAND3X1_211 ( );
FILL FILL_4_NAND3X1_211 ( );
FILL FILL_5_NAND3X1_211 ( );
FILL FILL_6_NAND3X1_211 ( );
FILL FILL_7_NAND3X1_211 ( );
FILL FILL_8_NAND3X1_211 ( );
FILL FILL_9_NAND3X1_211 ( );
FILL FILL_0_OAI21X1_37 ( );
FILL FILL_1_OAI21X1_37 ( );
FILL FILL_2_OAI21X1_37 ( );
FILL FILL_3_OAI21X1_37 ( );
FILL FILL_4_OAI21X1_37 ( );
FILL FILL_5_OAI21X1_37 ( );
FILL FILL_6_OAI21X1_37 ( );
FILL FILL_7_OAI21X1_37 ( );
FILL FILL_8_OAI21X1_37 ( );
FILL FILL_9_OAI21X1_37 ( );
FILL FILL_0_INVX1_152 ( );
FILL FILL_1_INVX1_152 ( );
FILL FILL_2_INVX1_152 ( );
FILL FILL_3_INVX1_152 ( );
FILL FILL_4_INVX1_152 ( );
FILL FILL_0_AOI21X1_15 ( );
FILL FILL_1_AOI21X1_15 ( );
FILL FILL_2_AOI21X1_15 ( );
FILL FILL_3_AOI21X1_15 ( );
FILL FILL_4_AOI21X1_15 ( );
FILL FILL_5_AOI21X1_15 ( );
FILL FILL_6_AOI21X1_15 ( );
FILL FILL_7_AOI21X1_15 ( );
FILL FILL_8_AOI21X1_15 ( );
FILL FILL_9_AOI21X1_15 ( );
FILL FILL_0_NAND3X1_145 ( );
FILL FILL_1_NAND3X1_145 ( );
FILL FILL_2_NAND3X1_145 ( );
FILL FILL_3_NAND3X1_145 ( );
FILL FILL_4_NAND3X1_145 ( );
FILL FILL_5_NAND3X1_145 ( );
FILL FILL_6_NAND3X1_145 ( );
FILL FILL_7_NAND3X1_145 ( );
FILL FILL_8_NAND3X1_145 ( );
FILL FILL_0_NAND3X1_151 ( );
FILL FILL_1_NAND3X1_151 ( );
FILL FILL_2_NAND3X1_151 ( );
FILL FILL_3_NAND3X1_151 ( );
FILL FILL_4_NAND3X1_151 ( );
FILL FILL_5_NAND3X1_151 ( );
FILL FILL_6_NAND3X1_151 ( );
FILL FILL_7_NAND3X1_151 ( );
FILL FILL_8_NAND3X1_151 ( );
FILL FILL_9_NAND3X1_151 ( );
FILL FILL_0_OAI21X1_30 ( );
FILL FILL_1_OAI21X1_30 ( );
FILL FILL_2_OAI21X1_30 ( );
FILL FILL_3_OAI21X1_30 ( );
FILL FILL_4_OAI21X1_30 ( );
FILL FILL_5_OAI21X1_30 ( );
FILL FILL_6_OAI21X1_30 ( );
FILL FILL_7_OAI21X1_30 ( );
FILL FILL_8_OAI21X1_30 ( );
FILL FILL_9_OAI21X1_30 ( );
FILL FILL_0_INVX1_138 ( );
FILL FILL_1_INVX1_138 ( );
FILL FILL_2_INVX1_138 ( );
FILL FILL_3_INVX1_138 ( );
FILL FILL_4_INVX1_138 ( );
FILL FILL_0_INVX1_139 ( );
FILL FILL_1_INVX1_139 ( );
FILL FILL_2_INVX1_139 ( );
FILL FILL_3_INVX1_139 ( );
FILL FILL_4_INVX1_139 ( );
FILL FILL_0_DFFPOSX1_22 ( );
FILL FILL_1_DFFPOSX1_22 ( );
FILL FILL_2_DFFPOSX1_22 ( );
FILL FILL_3_DFFPOSX1_22 ( );
FILL FILL_4_DFFPOSX1_22 ( );
FILL FILL_5_DFFPOSX1_22 ( );
FILL FILL_6_DFFPOSX1_22 ( );
FILL FILL_7_DFFPOSX1_22 ( );
FILL FILL_8_DFFPOSX1_22 ( );
FILL FILL_9_DFFPOSX1_22 ( );
FILL FILL_10_DFFPOSX1_22 ( );
FILL FILL_11_DFFPOSX1_22 ( );
FILL FILL_12_DFFPOSX1_22 ( );
FILL FILL_13_DFFPOSX1_22 ( );
FILL FILL_14_DFFPOSX1_22 ( );
FILL FILL_15_DFFPOSX1_22 ( );
FILL FILL_16_DFFPOSX1_22 ( );
FILL FILL_17_DFFPOSX1_22 ( );
FILL FILL_18_DFFPOSX1_22 ( );
FILL FILL_19_DFFPOSX1_22 ( );
FILL FILL_20_DFFPOSX1_22 ( );
FILL FILL_21_DFFPOSX1_22 ( );
FILL FILL_22_DFFPOSX1_22 ( );
FILL FILL_23_DFFPOSX1_22 ( );
FILL FILL_24_DFFPOSX1_22 ( );
FILL FILL_25_DFFPOSX1_22 ( );
FILL FILL_26_DFFPOSX1_22 ( );
FILL FILL_27_DFFPOSX1_22 ( );
FILL FILL_0_INVX1_196 ( );
FILL FILL_1_INVX1_196 ( );
FILL FILL_2_INVX1_196 ( );
FILL FILL_3_INVX1_196 ( );
FILL FILL_0_CLKBUF1_44 ( );
FILL FILL_1_CLKBUF1_44 ( );
FILL FILL_2_CLKBUF1_44 ( );
FILL FILL_3_CLKBUF1_44 ( );
FILL FILL_4_CLKBUF1_44 ( );
FILL FILL_5_CLKBUF1_44 ( );
FILL FILL_6_CLKBUF1_44 ( );
FILL FILL_7_CLKBUF1_44 ( );
FILL FILL_8_CLKBUF1_44 ( );
FILL FILL_9_CLKBUF1_44 ( );
FILL FILL_10_CLKBUF1_44 ( );
FILL FILL_11_CLKBUF1_44 ( );
FILL FILL_12_CLKBUF1_44 ( );
FILL FILL_13_CLKBUF1_44 ( );
FILL FILL_14_CLKBUF1_44 ( );
FILL FILL_15_CLKBUF1_44 ( );
FILL FILL_16_CLKBUF1_44 ( );
FILL FILL_17_CLKBUF1_44 ( );
FILL FILL_18_CLKBUF1_44 ( );
FILL FILL_19_CLKBUF1_44 ( );
FILL FILL_20_CLKBUF1_44 ( );
FILL FILL_0_NAND2X1_151 ( );
FILL FILL_1_NAND2X1_151 ( );
FILL FILL_2_NAND2X1_151 ( );
FILL FILL_3_NAND2X1_151 ( );
FILL FILL_4_NAND2X1_151 ( );
FILL FILL_5_NAND2X1_151 ( );
FILL FILL_6_NAND2X1_151 ( );
FILL FILL_0_AOI21X1_51 ( );
FILL FILL_1_AOI21X1_51 ( );
FILL FILL_2_AOI21X1_51 ( );
FILL FILL_3_AOI21X1_51 ( );
FILL FILL_4_AOI21X1_51 ( );
FILL FILL_5_AOI21X1_51 ( );
FILL FILL_6_AOI21X1_51 ( );
FILL FILL_7_AOI21X1_51 ( );
FILL FILL_8_AOI21X1_51 ( );
FILL FILL_0_NAND3X1_136 ( );
FILL FILL_1_NAND3X1_136 ( );
FILL FILL_2_NAND3X1_136 ( );
FILL FILL_3_NAND3X1_136 ( );
FILL FILL_4_NAND3X1_136 ( );
FILL FILL_5_NAND3X1_136 ( );
FILL FILL_6_NAND3X1_136 ( );
FILL FILL_7_NAND3X1_136 ( );
FILL FILL_8_NAND3X1_136 ( );
FILL FILL_0_AOI21X1_6 ( );
FILL FILL_1_AOI21X1_6 ( );
FILL FILL_2_AOI21X1_6 ( );
FILL FILL_3_AOI21X1_6 ( );
FILL FILL_4_AOI21X1_6 ( );
FILL FILL_5_AOI21X1_6 ( );
FILL FILL_6_AOI21X1_6 ( );
FILL FILL_7_AOI21X1_6 ( );
FILL FILL_8_AOI21X1_6 ( );
FILL FILL_9_AOI21X1_6 ( );
FILL FILL_0_CLKBUF1_32 ( );
FILL FILL_1_CLKBUF1_32 ( );
FILL FILL_2_CLKBUF1_32 ( );
FILL FILL_3_CLKBUF1_32 ( );
FILL FILL_4_CLKBUF1_32 ( );
FILL FILL_5_CLKBUF1_32 ( );
FILL FILL_6_CLKBUF1_32 ( );
FILL FILL_7_CLKBUF1_32 ( );
FILL FILL_8_CLKBUF1_32 ( );
FILL FILL_9_CLKBUF1_32 ( );
FILL FILL_10_CLKBUF1_32 ( );
FILL FILL_11_CLKBUF1_32 ( );
FILL FILL_12_CLKBUF1_32 ( );
FILL FILL_13_CLKBUF1_32 ( );
FILL FILL_14_CLKBUF1_32 ( );
FILL FILL_15_CLKBUF1_32 ( );
FILL FILL_16_CLKBUF1_32 ( );
FILL FILL_17_CLKBUF1_32 ( );
FILL FILL_18_CLKBUF1_32 ( );
FILL FILL_19_CLKBUF1_32 ( );
FILL FILL_20_CLKBUF1_32 ( );
FILL FILL_0_AND2X2_41 ( );
FILL FILL_1_AND2X2_41 ( );
FILL FILL_2_AND2X2_41 ( );
FILL FILL_3_AND2X2_41 ( );
FILL FILL_4_AND2X2_41 ( );
FILL FILL_5_AND2X2_41 ( );
FILL FILL_6_AND2X2_41 ( );
FILL FILL_7_AND2X2_41 ( );
FILL FILL_8_AND2X2_41 ( );
FILL FILL_0_DFFSR_81 ( );
FILL FILL_1_DFFSR_81 ( );
FILL FILL_2_DFFSR_81 ( );
FILL FILL_3_DFFSR_81 ( );
FILL FILL_4_DFFSR_81 ( );
FILL FILL_5_DFFSR_81 ( );
FILL FILL_6_DFFSR_81 ( );
FILL FILL_7_DFFSR_81 ( );
FILL FILL_8_DFFSR_81 ( );
FILL FILL_9_DFFSR_81 ( );
FILL FILL_10_DFFSR_81 ( );
FILL FILL_11_DFFSR_81 ( );
FILL FILL_12_DFFSR_81 ( );
FILL FILL_13_DFFSR_81 ( );
FILL FILL_14_DFFSR_81 ( );
FILL FILL_15_DFFSR_81 ( );
FILL FILL_16_DFFSR_81 ( );
FILL FILL_17_DFFSR_81 ( );
FILL FILL_18_DFFSR_81 ( );
FILL FILL_19_DFFSR_81 ( );
FILL FILL_20_DFFSR_81 ( );
FILL FILL_21_DFFSR_81 ( );
FILL FILL_22_DFFSR_81 ( );
FILL FILL_23_DFFSR_81 ( );
FILL FILL_24_DFFSR_81 ( );
FILL FILL_25_DFFSR_81 ( );
FILL FILL_26_DFFSR_81 ( );
FILL FILL_27_DFFSR_81 ( );
FILL FILL_28_DFFSR_81 ( );
FILL FILL_29_DFFSR_81 ( );
FILL FILL_30_DFFSR_81 ( );
FILL FILL_31_DFFSR_81 ( );
FILL FILL_32_DFFSR_81 ( );
FILL FILL_33_DFFSR_81 ( );
FILL FILL_34_DFFSR_81 ( );
FILL FILL_35_DFFSR_81 ( );
FILL FILL_36_DFFSR_81 ( );
FILL FILL_37_DFFSR_81 ( );
FILL FILL_38_DFFSR_81 ( );
FILL FILL_39_DFFSR_81 ( );
FILL FILL_40_DFFSR_81 ( );
FILL FILL_41_DFFSR_81 ( );
FILL FILL_42_DFFSR_81 ( );
FILL FILL_43_DFFSR_81 ( );
FILL FILL_44_DFFSR_81 ( );
FILL FILL_45_DFFSR_81 ( );
FILL FILL_46_DFFSR_81 ( );
FILL FILL_47_DFFSR_81 ( );
FILL FILL_48_DFFSR_81 ( );
FILL FILL_49_DFFSR_81 ( );
FILL FILL_50_DFFSR_81 ( );
FILL FILL_51_DFFSR_81 ( );
FILL FILL_0_DFFSR_244 ( );
FILL FILL_1_DFFSR_244 ( );
FILL FILL_2_DFFSR_244 ( );
FILL FILL_3_DFFSR_244 ( );
FILL FILL_4_DFFSR_244 ( );
FILL FILL_5_DFFSR_244 ( );
FILL FILL_6_DFFSR_244 ( );
FILL FILL_7_DFFSR_244 ( );
FILL FILL_8_DFFSR_244 ( );
FILL FILL_9_DFFSR_244 ( );
FILL FILL_10_DFFSR_244 ( );
FILL FILL_11_DFFSR_244 ( );
FILL FILL_12_DFFSR_244 ( );
FILL FILL_13_DFFSR_244 ( );
FILL FILL_14_DFFSR_244 ( );
FILL FILL_15_DFFSR_244 ( );
FILL FILL_16_DFFSR_244 ( );
FILL FILL_17_DFFSR_244 ( );
FILL FILL_18_DFFSR_244 ( );
FILL FILL_19_DFFSR_244 ( );
FILL FILL_20_DFFSR_244 ( );
FILL FILL_21_DFFSR_244 ( );
FILL FILL_22_DFFSR_244 ( );
FILL FILL_23_DFFSR_244 ( );
FILL FILL_24_DFFSR_244 ( );
FILL FILL_25_DFFSR_244 ( );
FILL FILL_26_DFFSR_244 ( );
FILL FILL_27_DFFSR_244 ( );
FILL FILL_28_DFFSR_244 ( );
FILL FILL_29_DFFSR_244 ( );
FILL FILL_30_DFFSR_244 ( );
FILL FILL_31_DFFSR_244 ( );
FILL FILL_32_DFFSR_244 ( );
FILL FILL_33_DFFSR_244 ( );
FILL FILL_34_DFFSR_244 ( );
FILL FILL_35_DFFSR_244 ( );
FILL FILL_36_DFFSR_244 ( );
FILL FILL_37_DFFSR_244 ( );
FILL FILL_38_DFFSR_244 ( );
FILL FILL_39_DFFSR_244 ( );
FILL FILL_40_DFFSR_244 ( );
FILL FILL_41_DFFSR_244 ( );
FILL FILL_42_DFFSR_244 ( );
FILL FILL_43_DFFSR_244 ( );
FILL FILL_44_DFFSR_244 ( );
FILL FILL_45_DFFSR_244 ( );
FILL FILL_46_DFFSR_244 ( );
FILL FILL_47_DFFSR_244 ( );
FILL FILL_48_DFFSR_244 ( );
FILL FILL_49_DFFSR_244 ( );
FILL FILL_50_DFFSR_244 ( );
FILL FILL_0_NAND3X1_88 ( );
FILL FILL_1_NAND3X1_88 ( );
FILL FILL_2_NAND3X1_88 ( );
FILL FILL_3_NAND3X1_88 ( );
FILL FILL_4_NAND3X1_88 ( );
FILL FILL_5_NAND3X1_88 ( );
FILL FILL_6_NAND3X1_88 ( );
FILL FILL_7_NAND3X1_88 ( );
FILL FILL_8_NAND3X1_88 ( );
FILL FILL_9_NAND3X1_88 ( );
FILL FILL_0_NOR2X1_41 ( );
FILL FILL_1_NOR2X1_41 ( );
FILL FILL_2_NOR2X1_41 ( );
FILL FILL_3_NOR2X1_41 ( );
FILL FILL_4_NOR2X1_41 ( );
FILL FILL_5_NOR2X1_41 ( );
FILL FILL_6_NOR2X1_41 ( );
FILL FILL_0_INVX1_80 ( );
FILL FILL_1_INVX1_80 ( );
FILL FILL_2_INVX1_80 ( );
FILL FILL_3_INVX1_80 ( );
FILL FILL_4_INVX1_80 ( );
FILL FILL_0_NAND3X1_105 ( );
FILL FILL_1_NAND3X1_105 ( );
FILL FILL_2_NAND3X1_105 ( );
FILL FILL_3_NAND3X1_105 ( );
FILL FILL_4_NAND3X1_105 ( );
FILL FILL_5_NAND3X1_105 ( );
FILL FILL_6_NAND3X1_105 ( );
FILL FILL_7_NAND3X1_105 ( );
FILL FILL_8_NAND3X1_105 ( );
FILL FILL_0_OAI22X1_31 ( );
FILL FILL_1_OAI22X1_31 ( );
FILL FILL_2_OAI22X1_31 ( );
FILL FILL_3_OAI22X1_31 ( );
FILL FILL_4_OAI22X1_31 ( );
FILL FILL_5_OAI22X1_31 ( );
FILL FILL_6_OAI22X1_31 ( );
FILL FILL_7_OAI22X1_31 ( );
FILL FILL_8_OAI22X1_31 ( );
FILL FILL_9_OAI22X1_31 ( );
FILL FILL_10_OAI22X1_31 ( );
FILL FILL_11_OAI22X1_31 ( );
FILL FILL_0_INVX1_77 ( );
FILL FILL_1_INVX1_77 ( );
FILL FILL_2_INVX1_77 ( );
FILL FILL_3_INVX1_77 ( );
FILL FILL_0_DFFSR_187 ( );
FILL FILL_1_DFFSR_187 ( );
FILL FILL_2_DFFSR_187 ( );
FILL FILL_3_DFFSR_187 ( );
FILL FILL_4_DFFSR_187 ( );
FILL FILL_5_DFFSR_187 ( );
FILL FILL_6_DFFSR_187 ( );
FILL FILL_7_DFFSR_187 ( );
FILL FILL_8_DFFSR_187 ( );
FILL FILL_9_DFFSR_187 ( );
FILL FILL_10_DFFSR_187 ( );
FILL FILL_11_DFFSR_187 ( );
FILL FILL_12_DFFSR_187 ( );
FILL FILL_13_DFFSR_187 ( );
FILL FILL_14_DFFSR_187 ( );
FILL FILL_15_DFFSR_187 ( );
FILL FILL_16_DFFSR_187 ( );
FILL FILL_17_DFFSR_187 ( );
FILL FILL_18_DFFSR_187 ( );
FILL FILL_19_DFFSR_187 ( );
FILL FILL_20_DFFSR_187 ( );
FILL FILL_21_DFFSR_187 ( );
FILL FILL_22_DFFSR_187 ( );
FILL FILL_23_DFFSR_187 ( );
FILL FILL_24_DFFSR_187 ( );
FILL FILL_25_DFFSR_187 ( );
FILL FILL_26_DFFSR_187 ( );
FILL FILL_27_DFFSR_187 ( );
FILL FILL_28_DFFSR_187 ( );
FILL FILL_29_DFFSR_187 ( );
FILL FILL_30_DFFSR_187 ( );
FILL FILL_31_DFFSR_187 ( );
FILL FILL_32_DFFSR_187 ( );
FILL FILL_33_DFFSR_187 ( );
FILL FILL_34_DFFSR_187 ( );
FILL FILL_35_DFFSR_187 ( );
FILL FILL_36_DFFSR_187 ( );
FILL FILL_37_DFFSR_187 ( );
FILL FILL_38_DFFSR_187 ( );
FILL FILL_39_DFFSR_187 ( );
FILL FILL_40_DFFSR_187 ( );
FILL FILL_41_DFFSR_187 ( );
FILL FILL_42_DFFSR_187 ( );
FILL FILL_43_DFFSR_187 ( );
FILL FILL_44_DFFSR_187 ( );
FILL FILL_45_DFFSR_187 ( );
FILL FILL_46_DFFSR_187 ( );
FILL FILL_47_DFFSR_187 ( );
FILL FILL_48_DFFSR_187 ( );
FILL FILL_49_DFFSR_187 ( );
FILL FILL_50_DFFSR_187 ( );
FILL FILL_0_OAI22X1_44 ( );
FILL FILL_1_OAI22X1_44 ( );
FILL FILL_2_OAI22X1_44 ( );
FILL FILL_3_OAI22X1_44 ( );
FILL FILL_4_OAI22X1_44 ( );
FILL FILL_5_OAI22X1_44 ( );
FILL FILL_6_OAI22X1_44 ( );
FILL FILL_7_OAI22X1_44 ( );
FILL FILL_8_OAI22X1_44 ( );
FILL FILL_9_OAI22X1_44 ( );
FILL FILL_10_OAI22X1_44 ( );
FILL FILL_11_OAI22X1_44 ( );
FILL FILL_0_NOR2X1_53 ( );
FILL FILL_1_NOR2X1_53 ( );
FILL FILL_2_NOR2X1_53 ( );
FILL FILL_3_NOR2X1_53 ( );
FILL FILL_4_NOR2X1_53 ( );
FILL FILL_5_NOR2X1_53 ( );
FILL FILL_6_NOR2X1_53 ( );
FILL FILL_0_BUFX2_66 ( );
FILL FILL_1_BUFX2_66 ( );
FILL FILL_2_BUFX2_66 ( );
FILL FILL_3_BUFX2_66 ( );
FILL FILL_4_BUFX2_66 ( );
FILL FILL_5_BUFX2_66 ( );
FILL FILL_6_BUFX2_66 ( );
FILL FILL_0_DFFSR_194 ( );
FILL FILL_1_DFFSR_194 ( );
FILL FILL_2_DFFSR_194 ( );
FILL FILL_3_DFFSR_194 ( );
FILL FILL_4_DFFSR_194 ( );
FILL FILL_5_DFFSR_194 ( );
FILL FILL_6_DFFSR_194 ( );
FILL FILL_7_DFFSR_194 ( );
FILL FILL_8_DFFSR_194 ( );
FILL FILL_9_DFFSR_194 ( );
FILL FILL_10_DFFSR_194 ( );
FILL FILL_11_DFFSR_194 ( );
FILL FILL_12_DFFSR_194 ( );
FILL FILL_13_DFFSR_194 ( );
FILL FILL_14_DFFSR_194 ( );
FILL FILL_15_DFFSR_194 ( );
FILL FILL_16_DFFSR_194 ( );
FILL FILL_17_DFFSR_194 ( );
FILL FILL_18_DFFSR_194 ( );
FILL FILL_19_DFFSR_194 ( );
FILL FILL_20_DFFSR_194 ( );
FILL FILL_21_DFFSR_194 ( );
FILL FILL_22_DFFSR_194 ( );
FILL FILL_23_DFFSR_194 ( );
FILL FILL_24_DFFSR_194 ( );
FILL FILL_25_DFFSR_194 ( );
FILL FILL_26_DFFSR_194 ( );
FILL FILL_27_DFFSR_194 ( );
FILL FILL_28_DFFSR_194 ( );
FILL FILL_29_DFFSR_194 ( );
FILL FILL_30_DFFSR_194 ( );
FILL FILL_31_DFFSR_194 ( );
FILL FILL_32_DFFSR_194 ( );
FILL FILL_33_DFFSR_194 ( );
FILL FILL_34_DFFSR_194 ( );
FILL FILL_35_DFFSR_194 ( );
FILL FILL_36_DFFSR_194 ( );
FILL FILL_37_DFFSR_194 ( );
FILL FILL_38_DFFSR_194 ( );
FILL FILL_39_DFFSR_194 ( );
FILL FILL_40_DFFSR_194 ( );
FILL FILL_41_DFFSR_194 ( );
FILL FILL_42_DFFSR_194 ( );
FILL FILL_43_DFFSR_194 ( );
FILL FILL_44_DFFSR_194 ( );
FILL FILL_45_DFFSR_194 ( );
FILL FILL_46_DFFSR_194 ( );
FILL FILL_47_DFFSR_194 ( );
FILL FILL_48_DFFSR_194 ( );
FILL FILL_49_DFFSR_194 ( );
FILL FILL_50_DFFSR_194 ( );
FILL FILL_51_DFFSR_194 ( );
FILL FILL_0_OAI21X1_48 ( );
FILL FILL_1_OAI21X1_48 ( );
FILL FILL_2_OAI21X1_48 ( );
FILL FILL_3_OAI21X1_48 ( );
FILL FILL_4_OAI21X1_48 ( );
FILL FILL_5_OAI21X1_48 ( );
FILL FILL_6_OAI21X1_48 ( );
FILL FILL_7_OAI21X1_48 ( );
FILL FILL_8_OAI21X1_48 ( );
FILL FILL_0_INVX1_150 ( );
FILL FILL_1_INVX1_150 ( );
FILL FILL_2_INVX1_150 ( );
FILL FILL_3_INVX1_150 ( );
FILL FILL_4_INVX1_150 ( );
FILL FILL_0_INVX1_164 ( );
FILL FILL_1_INVX1_164 ( );
FILL FILL_2_INVX1_164 ( );
FILL FILL_3_INVX1_164 ( );
FILL FILL_4_INVX1_164 ( );
FILL FILL_0_NAND3X1_210 ( );
FILL FILL_1_NAND3X1_210 ( );
FILL FILL_2_NAND3X1_210 ( );
FILL FILL_3_NAND3X1_210 ( );
FILL FILL_4_NAND3X1_210 ( );
FILL FILL_5_NAND3X1_210 ( );
FILL FILL_6_NAND3X1_210 ( );
FILL FILL_7_NAND3X1_210 ( );
FILL FILL_8_NAND3X1_210 ( );
FILL FILL_0_NAND3X1_206 ( );
FILL FILL_1_NAND3X1_206 ( );
FILL FILL_2_NAND3X1_206 ( );
FILL FILL_3_NAND3X1_206 ( );
FILL FILL_4_NAND3X1_206 ( );
FILL FILL_5_NAND3X1_206 ( );
FILL FILL_6_NAND3X1_206 ( );
FILL FILL_7_NAND3X1_206 ( );
FILL FILL_8_NAND3X1_206 ( );
FILL FILL_0_AOI21X1_10 ( );
FILL FILL_1_AOI21X1_10 ( );
FILL FILL_2_AOI21X1_10 ( );
FILL FILL_3_AOI21X1_10 ( );
FILL FILL_4_AOI21X1_10 ( );
FILL FILL_5_AOI21X1_10 ( );
FILL FILL_6_AOI21X1_10 ( );
FILL FILL_7_AOI21X1_10 ( );
FILL FILL_8_AOI21X1_10 ( );
FILL FILL_0_INVX1_143 ( );
FILL FILL_1_INVX1_143 ( );
FILL FILL_2_INVX1_143 ( );
FILL FILL_3_INVX1_143 ( );
FILL FILL_0_NAND2X1_66 ( );
FILL FILL_1_NAND2X1_66 ( );
FILL FILL_2_NAND2X1_66 ( );
FILL FILL_3_NAND2X1_66 ( );
FILL FILL_4_NAND2X1_66 ( );
FILL FILL_5_NAND2X1_66 ( );
FILL FILL_6_NAND2X1_66 ( );
FILL FILL_0_NAND3X1_148 ( );
FILL FILL_1_NAND3X1_148 ( );
FILL FILL_2_NAND3X1_148 ( );
FILL FILL_3_NAND3X1_148 ( );
FILL FILL_4_NAND3X1_148 ( );
FILL FILL_5_NAND3X1_148 ( );
FILL FILL_6_NAND3X1_148 ( );
FILL FILL_7_NAND3X1_148 ( );
FILL FILL_8_NAND3X1_148 ( );
FILL FILL_9_NAND3X1_148 ( );
FILL FILL_0_AOI21X1_14 ( );
FILL FILL_1_AOI21X1_14 ( );
FILL FILL_2_AOI21X1_14 ( );
FILL FILL_3_AOI21X1_14 ( );
FILL FILL_4_AOI21X1_14 ( );
FILL FILL_5_AOI21X1_14 ( );
FILL FILL_6_AOI21X1_14 ( );
FILL FILL_7_AOI21X1_14 ( );
FILL FILL_8_AOI21X1_14 ( );
FILL FILL_0_NAND2X1_62 ( );
FILL FILL_1_NAND2X1_62 ( );
FILL FILL_2_NAND2X1_62 ( );
FILL FILL_3_NAND2X1_62 ( );
FILL FILL_4_NAND2X1_62 ( );
FILL FILL_5_NAND2X1_62 ( );
FILL FILL_6_NAND2X1_62 ( );
FILL FILL_0_NAND2X1_58 ( );
FILL FILL_1_NAND2X1_58 ( );
FILL FILL_2_NAND2X1_58 ( );
FILL FILL_3_NAND2X1_58 ( );
FILL FILL_4_NAND2X1_58 ( );
FILL FILL_5_NAND2X1_58 ( );
FILL FILL_6_NAND2X1_58 ( );
FILL FILL_0_BUFX2_58 ( );
FILL FILL_1_BUFX2_58 ( );
FILL FILL_2_BUFX2_58 ( );
FILL FILL_3_BUFX2_58 ( );
FILL FILL_4_BUFX2_58 ( );
FILL FILL_5_BUFX2_58 ( );
FILL FILL_6_BUFX2_58 ( );
FILL FILL_0_DFFSR_271 ( );
FILL FILL_1_DFFSR_271 ( );
FILL FILL_2_DFFSR_271 ( );
FILL FILL_3_DFFSR_271 ( );
FILL FILL_4_DFFSR_271 ( );
FILL FILL_5_DFFSR_271 ( );
FILL FILL_6_DFFSR_271 ( );
FILL FILL_7_DFFSR_271 ( );
FILL FILL_8_DFFSR_271 ( );
FILL FILL_9_DFFSR_271 ( );
FILL FILL_10_DFFSR_271 ( );
FILL FILL_11_DFFSR_271 ( );
FILL FILL_12_DFFSR_271 ( );
FILL FILL_13_DFFSR_271 ( );
FILL FILL_14_DFFSR_271 ( );
FILL FILL_15_DFFSR_271 ( );
FILL FILL_16_DFFSR_271 ( );
FILL FILL_17_DFFSR_271 ( );
FILL FILL_18_DFFSR_271 ( );
FILL FILL_19_DFFSR_271 ( );
FILL FILL_20_DFFSR_271 ( );
FILL FILL_21_DFFSR_271 ( );
FILL FILL_22_DFFSR_271 ( );
FILL FILL_23_DFFSR_271 ( );
FILL FILL_24_DFFSR_271 ( );
FILL FILL_25_DFFSR_271 ( );
FILL FILL_26_DFFSR_271 ( );
FILL FILL_27_DFFSR_271 ( );
FILL FILL_28_DFFSR_271 ( );
FILL FILL_29_DFFSR_271 ( );
FILL FILL_30_DFFSR_271 ( );
FILL FILL_31_DFFSR_271 ( );
FILL FILL_32_DFFSR_271 ( );
FILL FILL_33_DFFSR_271 ( );
FILL FILL_34_DFFSR_271 ( );
FILL FILL_35_DFFSR_271 ( );
FILL FILL_36_DFFSR_271 ( );
FILL FILL_37_DFFSR_271 ( );
FILL FILL_38_DFFSR_271 ( );
FILL FILL_39_DFFSR_271 ( );
FILL FILL_40_DFFSR_271 ( );
FILL FILL_41_DFFSR_271 ( );
FILL FILL_42_DFFSR_271 ( );
FILL FILL_43_DFFSR_271 ( );
FILL FILL_44_DFFSR_271 ( );
FILL FILL_45_DFFSR_271 ( );
FILL FILL_46_DFFSR_271 ( );
FILL FILL_47_DFFSR_271 ( );
FILL FILL_48_DFFSR_271 ( );
FILL FILL_49_DFFSR_271 ( );
FILL FILL_50_DFFSR_271 ( );
FILL FILL_51_DFFSR_271 ( );
FILL FILL_0_NAND2X1_166 ( );
FILL FILL_1_NAND2X1_166 ( );
FILL FILL_2_NAND2X1_166 ( );
FILL FILL_3_NAND2X1_166 ( );
FILL FILL_4_NAND2X1_166 ( );
FILL FILL_5_NAND2X1_166 ( );
FILL FILL_6_NAND2X1_166 ( );
FILL FILL_0_NAND3X1_135 ( );
FILL FILL_1_NAND3X1_135 ( );
FILL FILL_2_NAND3X1_135 ( );
FILL FILL_3_NAND3X1_135 ( );
FILL FILL_4_NAND3X1_135 ( );
FILL FILL_5_NAND3X1_135 ( );
FILL FILL_6_NAND3X1_135 ( );
FILL FILL_7_NAND3X1_135 ( );
FILL FILL_8_NAND3X1_135 ( );
FILL FILL_0_CLKBUF1_49 ( );
FILL FILL_1_CLKBUF1_49 ( );
FILL FILL_2_CLKBUF1_49 ( );
FILL FILL_3_CLKBUF1_49 ( );
FILL FILL_4_CLKBUF1_49 ( );
FILL FILL_5_CLKBUF1_49 ( );
FILL FILL_6_CLKBUF1_49 ( );
FILL FILL_7_CLKBUF1_49 ( );
FILL FILL_8_CLKBUF1_49 ( );
FILL FILL_9_CLKBUF1_49 ( );
FILL FILL_10_CLKBUF1_49 ( );
FILL FILL_11_CLKBUF1_49 ( );
FILL FILL_12_CLKBUF1_49 ( );
FILL FILL_13_CLKBUF1_49 ( );
FILL FILL_14_CLKBUF1_49 ( );
FILL FILL_15_CLKBUF1_49 ( );
FILL FILL_16_CLKBUF1_49 ( );
FILL FILL_17_CLKBUF1_49 ( );
FILL FILL_18_CLKBUF1_49 ( );
FILL FILL_19_CLKBUF1_49 ( );
FILL FILL_20_CLKBUF1_49 ( );
FILL FILL_0_DFFPOSX1_13 ( );
FILL FILL_1_DFFPOSX1_13 ( );
FILL FILL_2_DFFPOSX1_13 ( );
FILL FILL_3_DFFPOSX1_13 ( );
FILL FILL_4_DFFPOSX1_13 ( );
FILL FILL_5_DFFPOSX1_13 ( );
FILL FILL_6_DFFPOSX1_13 ( );
FILL FILL_7_DFFPOSX1_13 ( );
FILL FILL_8_DFFPOSX1_13 ( );
FILL FILL_9_DFFPOSX1_13 ( );
FILL FILL_10_DFFPOSX1_13 ( );
FILL FILL_11_DFFPOSX1_13 ( );
FILL FILL_12_DFFPOSX1_13 ( );
FILL FILL_13_DFFPOSX1_13 ( );
FILL FILL_14_DFFPOSX1_13 ( );
FILL FILL_15_DFFPOSX1_13 ( );
FILL FILL_16_DFFPOSX1_13 ( );
FILL FILL_17_DFFPOSX1_13 ( );
FILL FILL_18_DFFPOSX1_13 ( );
FILL FILL_19_DFFPOSX1_13 ( );
FILL FILL_20_DFFPOSX1_13 ( );
FILL FILL_21_DFFPOSX1_13 ( );
FILL FILL_22_DFFPOSX1_13 ( );
FILL FILL_23_DFFPOSX1_13 ( );
FILL FILL_24_DFFPOSX1_13 ( );
FILL FILL_25_DFFPOSX1_13 ( );
FILL FILL_26_DFFPOSX1_13 ( );
FILL FILL_27_DFFPOSX1_13 ( );
FILL FILL_0_INVX1_213 ( );
FILL FILL_1_INVX1_213 ( );
FILL FILL_2_INVX1_213 ( );
FILL FILL_3_INVX1_213 ( );
FILL FILL_4_INVX1_213 ( );
FILL FILL_0_OR2X2_5 ( );
FILL FILL_1_OR2X2_5 ( );
FILL FILL_2_OR2X2_5 ( );
FILL FILL_3_OR2X2_5 ( );
FILL FILL_4_OR2X2_5 ( );
FILL FILL_5_OR2X2_5 ( );
FILL FILL_6_OR2X2_5 ( );
FILL FILL_7_OR2X2_5 ( );
FILL FILL_8_OR2X2_5 ( );
FILL FILL_0_OAI21X1_112 ( );
FILL FILL_1_OAI21X1_112 ( );
FILL FILL_2_OAI21X1_112 ( );
FILL FILL_3_OAI21X1_112 ( );
FILL FILL_4_OAI21X1_112 ( );
FILL FILL_5_OAI21X1_112 ( );
FILL FILL_6_OAI21X1_112 ( );
FILL FILL_7_OAI21X1_112 ( );
FILL FILL_8_OAI21X1_112 ( );
FILL FILL_9_OAI21X1_112 ( );
FILL FILL_0_INVX1_211 ( );
FILL FILL_1_INVX1_211 ( );
FILL FILL_2_INVX1_211 ( );
FILL FILL_3_INVX1_211 ( );
FILL FILL_4_INVX1_211 ( );
FILL FILL_0_BUFX2_3 ( );
FILL FILL_1_BUFX2_3 ( );
FILL FILL_2_BUFX2_3 ( );
FILL FILL_3_BUFX2_3 ( );
FILL FILL_4_BUFX2_3 ( );
FILL FILL_5_BUFX2_3 ( );
FILL FILL_6_BUFX2_3 ( );
FILL FILL_0_CLKBUF1_19 ( );
FILL FILL_1_CLKBUF1_19 ( );
FILL FILL_2_CLKBUF1_19 ( );
FILL FILL_3_CLKBUF1_19 ( );
FILL FILL_4_CLKBUF1_19 ( );
FILL FILL_5_CLKBUF1_19 ( );
FILL FILL_6_CLKBUF1_19 ( );
FILL FILL_7_CLKBUF1_19 ( );
FILL FILL_8_CLKBUF1_19 ( );
FILL FILL_9_CLKBUF1_19 ( );
FILL FILL_10_CLKBUF1_19 ( );
FILL FILL_11_CLKBUF1_19 ( );
FILL FILL_12_CLKBUF1_19 ( );
FILL FILL_13_CLKBUF1_19 ( );
FILL FILL_14_CLKBUF1_19 ( );
FILL FILL_15_CLKBUF1_19 ( );
FILL FILL_16_CLKBUF1_19 ( );
FILL FILL_17_CLKBUF1_19 ( );
FILL FILL_18_CLKBUF1_19 ( );
FILL FILL_19_CLKBUF1_19 ( );
FILL FILL_20_CLKBUF1_19 ( );
FILL FILL_0_INVX1_5 ( );
FILL FILL_1_INVX1_5 ( );
FILL FILL_2_INVX1_5 ( );
FILL FILL_3_INVX1_5 ( );
FILL FILL_4_INVX1_5 ( );
FILL FILL_0_INVX1_6 ( );
FILL FILL_1_INVX1_6 ( );
FILL FILL_2_INVX1_6 ( );
FILL FILL_3_INVX1_6 ( );
FILL FILL_4_INVX1_6 ( );
FILL FILL_0_INVX1_128 ( );
FILL FILL_1_INVX1_128 ( );
FILL FILL_2_INVX1_128 ( );
FILL FILL_3_INVX1_128 ( );
FILL FILL_4_INVX1_128 ( );
FILL FILL_0_CLKBUF1_17 ( );
FILL FILL_1_CLKBUF1_17 ( );
FILL FILL_2_CLKBUF1_17 ( );
FILL FILL_3_CLKBUF1_17 ( );
FILL FILL_4_CLKBUF1_17 ( );
FILL FILL_5_CLKBUF1_17 ( );
FILL FILL_6_CLKBUF1_17 ( );
FILL FILL_7_CLKBUF1_17 ( );
FILL FILL_8_CLKBUF1_17 ( );
FILL FILL_9_CLKBUF1_17 ( );
FILL FILL_10_CLKBUF1_17 ( );
FILL FILL_11_CLKBUF1_17 ( );
FILL FILL_12_CLKBUF1_17 ( );
FILL FILL_13_CLKBUF1_17 ( );
FILL FILL_14_CLKBUF1_17 ( );
FILL FILL_15_CLKBUF1_17 ( );
FILL FILL_16_CLKBUF1_17 ( );
FILL FILL_17_CLKBUF1_17 ( );
FILL FILL_18_CLKBUF1_17 ( );
FILL FILL_19_CLKBUF1_17 ( );
FILL FILL_20_CLKBUF1_17 ( );
FILL FILL_0_NAND2X1_43 ( );
FILL FILL_1_NAND2X1_43 ( );
FILL FILL_2_NAND2X1_43 ( );
FILL FILL_3_NAND2X1_43 ( );
FILL FILL_4_NAND2X1_43 ( );
FILL FILL_5_NAND2X1_43 ( );
FILL FILL_6_NAND2X1_43 ( );
FILL FILL_0_NAND2X1_38 ( );
FILL FILL_1_NAND2X1_38 ( );
FILL FILL_2_NAND2X1_38 ( );
FILL FILL_3_NAND2X1_38 ( );
FILL FILL_4_NAND2X1_38 ( );
FILL FILL_5_NAND2X1_38 ( );
FILL FILL_6_NAND2X1_38 ( );
FILL FILL_0_NAND3X1_108 ( );
FILL FILL_1_NAND3X1_108 ( );
FILL FILL_2_NAND3X1_108 ( );
FILL FILL_3_NAND3X1_108 ( );
FILL FILL_4_NAND3X1_108 ( );
FILL FILL_5_NAND3X1_108 ( );
FILL FILL_6_NAND3X1_108 ( );
FILL FILL_7_NAND3X1_108 ( );
FILL FILL_8_NAND3X1_108 ( );
FILL FILL_9_NAND3X1_108 ( );
FILL FILL_0_NOR2X1_42 ( );
FILL FILL_1_NOR2X1_42 ( );
FILL FILL_2_NOR2X1_42 ( );
FILL FILL_3_NOR2X1_42 ( );
FILL FILL_4_NOR2X1_42 ( );
FILL FILL_5_NOR2X1_42 ( );
FILL FILL_6_NOR2X1_42 ( );
FILL FILL_0_NAND2X1_48 ( );
FILL FILL_1_NAND2X1_48 ( );
FILL FILL_2_NAND2X1_48 ( );
FILL FILL_3_NAND2X1_48 ( );
FILL FILL_4_NAND2X1_48 ( );
FILL FILL_5_NAND2X1_48 ( );
FILL FILL_6_NAND2X1_48 ( );
FILL FILL_0_NAND3X1_107 ( );
FILL FILL_1_NAND3X1_107 ( );
FILL FILL_2_NAND3X1_107 ( );
FILL FILL_3_NAND3X1_107 ( );
FILL FILL_4_NAND3X1_107 ( );
FILL FILL_5_NAND3X1_107 ( );
FILL FILL_6_NAND3X1_107 ( );
FILL FILL_7_NAND3X1_107 ( );
FILL FILL_8_NAND3X1_107 ( );
FILL FILL_0_BUFX2_95 ( );
FILL FILL_1_BUFX2_95 ( );
FILL FILL_2_BUFX2_95 ( );
FILL FILL_3_BUFX2_95 ( );
FILL FILL_4_BUFX2_95 ( );
FILL FILL_5_BUFX2_95 ( );
FILL FILL_6_BUFX2_95 ( );
FILL FILL_0_BUFX2_25 ( );
FILL FILL_1_BUFX2_25 ( );
FILL FILL_2_BUFX2_25 ( );
FILL FILL_3_BUFX2_25 ( );
FILL FILL_4_BUFX2_25 ( );
FILL FILL_5_BUFX2_25 ( );
FILL FILL_6_BUFX2_25 ( );
FILL FILL_0_DFFSR_171 ( );
FILL FILL_1_DFFSR_171 ( );
FILL FILL_2_DFFSR_171 ( );
FILL FILL_3_DFFSR_171 ( );
FILL FILL_4_DFFSR_171 ( );
FILL FILL_5_DFFSR_171 ( );
FILL FILL_6_DFFSR_171 ( );
FILL FILL_7_DFFSR_171 ( );
FILL FILL_8_DFFSR_171 ( );
FILL FILL_9_DFFSR_171 ( );
FILL FILL_10_DFFSR_171 ( );
FILL FILL_11_DFFSR_171 ( );
FILL FILL_12_DFFSR_171 ( );
FILL FILL_13_DFFSR_171 ( );
FILL FILL_14_DFFSR_171 ( );
FILL FILL_15_DFFSR_171 ( );
FILL FILL_16_DFFSR_171 ( );
FILL FILL_17_DFFSR_171 ( );
FILL FILL_18_DFFSR_171 ( );
FILL FILL_19_DFFSR_171 ( );
FILL FILL_20_DFFSR_171 ( );
FILL FILL_21_DFFSR_171 ( );
FILL FILL_22_DFFSR_171 ( );
FILL FILL_23_DFFSR_171 ( );
FILL FILL_24_DFFSR_171 ( );
FILL FILL_25_DFFSR_171 ( );
FILL FILL_26_DFFSR_171 ( );
FILL FILL_27_DFFSR_171 ( );
FILL FILL_28_DFFSR_171 ( );
FILL FILL_29_DFFSR_171 ( );
FILL FILL_30_DFFSR_171 ( );
FILL FILL_31_DFFSR_171 ( );
FILL FILL_32_DFFSR_171 ( );
FILL FILL_33_DFFSR_171 ( );
FILL FILL_34_DFFSR_171 ( );
FILL FILL_35_DFFSR_171 ( );
FILL FILL_36_DFFSR_171 ( );
FILL FILL_37_DFFSR_171 ( );
FILL FILL_38_DFFSR_171 ( );
FILL FILL_39_DFFSR_171 ( );
FILL FILL_40_DFFSR_171 ( );
FILL FILL_41_DFFSR_171 ( );
FILL FILL_42_DFFSR_171 ( );
FILL FILL_43_DFFSR_171 ( );
FILL FILL_44_DFFSR_171 ( );
FILL FILL_45_DFFSR_171 ( );
FILL FILL_46_DFFSR_171 ( );
FILL FILL_47_DFFSR_171 ( );
FILL FILL_48_DFFSR_171 ( );
FILL FILL_49_DFFSR_171 ( );
FILL FILL_50_DFFSR_171 ( );
FILL FILL_0_OAI22X1_47 ( );
FILL FILL_1_OAI22X1_47 ( );
FILL FILL_2_OAI22X1_47 ( );
FILL FILL_3_OAI22X1_47 ( );
FILL FILL_4_OAI22X1_47 ( );
FILL FILL_5_OAI22X1_47 ( );
FILL FILL_6_OAI22X1_47 ( );
FILL FILL_7_OAI22X1_47 ( );
FILL FILL_8_OAI22X1_47 ( );
FILL FILL_9_OAI22X1_47 ( );
FILL FILL_10_OAI22X1_47 ( );
FILL FILL_0_DFFSR_138 ( );
FILL FILL_1_DFFSR_138 ( );
FILL FILL_2_DFFSR_138 ( );
FILL FILL_3_DFFSR_138 ( );
FILL FILL_4_DFFSR_138 ( );
FILL FILL_5_DFFSR_138 ( );
FILL FILL_6_DFFSR_138 ( );
FILL FILL_7_DFFSR_138 ( );
FILL FILL_8_DFFSR_138 ( );
FILL FILL_9_DFFSR_138 ( );
FILL FILL_10_DFFSR_138 ( );
FILL FILL_11_DFFSR_138 ( );
FILL FILL_12_DFFSR_138 ( );
FILL FILL_13_DFFSR_138 ( );
FILL FILL_14_DFFSR_138 ( );
FILL FILL_15_DFFSR_138 ( );
FILL FILL_16_DFFSR_138 ( );
FILL FILL_17_DFFSR_138 ( );
FILL FILL_18_DFFSR_138 ( );
FILL FILL_19_DFFSR_138 ( );
FILL FILL_20_DFFSR_138 ( );
FILL FILL_21_DFFSR_138 ( );
FILL FILL_22_DFFSR_138 ( );
FILL FILL_23_DFFSR_138 ( );
FILL FILL_24_DFFSR_138 ( );
FILL FILL_25_DFFSR_138 ( );
FILL FILL_26_DFFSR_138 ( );
FILL FILL_27_DFFSR_138 ( );
FILL FILL_28_DFFSR_138 ( );
FILL FILL_29_DFFSR_138 ( );
FILL FILL_30_DFFSR_138 ( );
FILL FILL_31_DFFSR_138 ( );
FILL FILL_32_DFFSR_138 ( );
FILL FILL_33_DFFSR_138 ( );
FILL FILL_34_DFFSR_138 ( );
FILL FILL_35_DFFSR_138 ( );
FILL FILL_36_DFFSR_138 ( );
FILL FILL_37_DFFSR_138 ( );
FILL FILL_38_DFFSR_138 ( );
FILL FILL_39_DFFSR_138 ( );
FILL FILL_40_DFFSR_138 ( );
FILL FILL_41_DFFSR_138 ( );
FILL FILL_42_DFFSR_138 ( );
FILL FILL_43_DFFSR_138 ( );
FILL FILL_44_DFFSR_138 ( );
FILL FILL_45_DFFSR_138 ( );
FILL FILL_46_DFFSR_138 ( );
FILL FILL_47_DFFSR_138 ( );
FILL FILL_48_DFFSR_138 ( );
FILL FILL_49_DFFSR_138 ( );
FILL FILL_50_DFFSR_138 ( );
FILL FILL_0_XNOR2X1_1 ( );
FILL FILL_1_XNOR2X1_1 ( );
FILL FILL_2_XNOR2X1_1 ( );
FILL FILL_3_XNOR2X1_1 ( );
FILL FILL_4_XNOR2X1_1 ( );
FILL FILL_5_XNOR2X1_1 ( );
FILL FILL_6_XNOR2X1_1 ( );
FILL FILL_7_XNOR2X1_1 ( );
FILL FILL_8_XNOR2X1_1 ( );
FILL FILL_9_XNOR2X1_1 ( );
FILL FILL_10_XNOR2X1_1 ( );
FILL FILL_11_XNOR2X1_1 ( );
FILL FILL_12_XNOR2X1_1 ( );
FILL FILL_13_XNOR2X1_1 ( );
FILL FILL_14_XNOR2X1_1 ( );
FILL FILL_15_XNOR2X1_1 ( );
FILL FILL_0_OAI21X1_36 ( );
FILL FILL_1_OAI21X1_36 ( );
FILL FILL_2_OAI21X1_36 ( );
FILL FILL_3_OAI21X1_36 ( );
FILL FILL_4_OAI21X1_36 ( );
FILL FILL_5_OAI21X1_36 ( );
FILL FILL_6_OAI21X1_36 ( );
FILL FILL_7_OAI21X1_36 ( );
FILL FILL_8_OAI21X1_36 ( );
FILL FILL_0_NAND3X1_184 ( );
FILL FILL_1_NAND3X1_184 ( );
FILL FILL_2_NAND3X1_184 ( );
FILL FILL_3_NAND3X1_184 ( );
FILL FILL_4_NAND3X1_184 ( );
FILL FILL_5_NAND3X1_184 ( );
FILL FILL_6_NAND3X1_184 ( );
FILL FILL_7_NAND3X1_184 ( );
FILL FILL_8_NAND3X1_184 ( );
FILL FILL_0_NAND3X1_162 ( );
FILL FILL_1_NAND3X1_162 ( );
FILL FILL_2_NAND3X1_162 ( );
FILL FILL_3_NAND3X1_162 ( );
FILL FILL_4_NAND3X1_162 ( );
FILL FILL_5_NAND3X1_162 ( );
FILL FILL_6_NAND3X1_162 ( );
FILL FILL_7_NAND3X1_162 ( );
FILL FILL_8_NAND3X1_162 ( );
FILL FILL_0_NAND3X1_159 ( );
FILL FILL_1_NAND3X1_159 ( );
FILL FILL_2_NAND3X1_159 ( );
FILL FILL_3_NAND3X1_159 ( );
FILL FILL_4_NAND3X1_159 ( );
FILL FILL_5_NAND3X1_159 ( );
FILL FILL_6_NAND3X1_159 ( );
FILL FILL_7_NAND3X1_159 ( );
FILL FILL_8_NAND3X1_159 ( );
FILL FILL_0_INVX1_135 ( );
FILL FILL_1_INVX1_135 ( );
FILL FILL_2_INVX1_135 ( );
FILL FILL_3_INVX1_135 ( );
FILL FILL_0_NAND3X1_146 ( );
FILL FILL_1_NAND3X1_146 ( );
FILL FILL_2_NAND3X1_146 ( );
FILL FILL_3_NAND3X1_146 ( );
FILL FILL_4_NAND3X1_146 ( );
FILL FILL_5_NAND3X1_146 ( );
FILL FILL_6_NAND3X1_146 ( );
FILL FILL_7_NAND3X1_146 ( );
FILL FILL_8_NAND3X1_146 ( );
FILL FILL_0_NAND3X1_143 ( );
FILL FILL_1_NAND3X1_143 ( );
FILL FILL_2_NAND3X1_143 ( );
FILL FILL_3_NAND3X1_143 ( );
FILL FILL_4_NAND3X1_143 ( );
FILL FILL_5_NAND3X1_143 ( );
FILL FILL_6_NAND3X1_143 ( );
FILL FILL_7_NAND3X1_143 ( );
FILL FILL_8_NAND3X1_143 ( );
FILL FILL_0_INVX1_144 ( );
FILL FILL_1_INVX1_144 ( );
FILL FILL_2_INVX1_144 ( );
FILL FILL_3_INVX1_144 ( );
FILL FILL_0_NAND3X1_139 ( );
FILL FILL_1_NAND3X1_139 ( );
FILL FILL_2_NAND3X1_139 ( );
FILL FILL_3_NAND3X1_139 ( );
FILL FILL_4_NAND3X1_139 ( );
FILL FILL_5_NAND3X1_139 ( );
FILL FILL_6_NAND3X1_139 ( );
FILL FILL_7_NAND3X1_139 ( );
FILL FILL_8_NAND3X1_139 ( );
FILL FILL_9_NAND3X1_139 ( );
FILL FILL_0_BUFX2_56 ( );
FILL FILL_1_BUFX2_56 ( );
FILL FILL_2_BUFX2_56 ( );
FILL FILL_3_BUFX2_56 ( );
FILL FILL_4_BUFX2_56 ( );
FILL FILL_5_BUFX2_56 ( );
FILL FILL_6_BUFX2_56 ( );
FILL FILL_0_INVX1_193 ( );
FILL FILL_1_INVX1_193 ( );
FILL FILL_2_INVX1_193 ( );
FILL FILL_3_INVX1_193 ( );
FILL FILL_0_DFFPOSX1_17 ( );
FILL FILL_1_DFFPOSX1_17 ( );
FILL FILL_2_DFFPOSX1_17 ( );
FILL FILL_3_DFFPOSX1_17 ( );
FILL FILL_4_DFFPOSX1_17 ( );
FILL FILL_5_DFFPOSX1_17 ( );
FILL FILL_6_DFFPOSX1_17 ( );
FILL FILL_7_DFFPOSX1_17 ( );
FILL FILL_8_DFFPOSX1_17 ( );
FILL FILL_9_DFFPOSX1_17 ( );
FILL FILL_10_DFFPOSX1_17 ( );
FILL FILL_11_DFFPOSX1_17 ( );
FILL FILL_12_DFFPOSX1_17 ( );
FILL FILL_13_DFFPOSX1_17 ( );
FILL FILL_14_DFFPOSX1_17 ( );
FILL FILL_15_DFFPOSX1_17 ( );
FILL FILL_16_DFFPOSX1_17 ( );
FILL FILL_17_DFFPOSX1_17 ( );
FILL FILL_18_DFFPOSX1_17 ( );
FILL FILL_19_DFFPOSX1_17 ( );
FILL FILL_20_DFFPOSX1_17 ( );
FILL FILL_21_DFFPOSX1_17 ( );
FILL FILL_22_DFFPOSX1_17 ( );
FILL FILL_23_DFFPOSX1_17 ( );
FILL FILL_24_DFFPOSX1_17 ( );
FILL FILL_25_DFFPOSX1_17 ( );
FILL FILL_26_DFFPOSX1_17 ( );
FILL FILL_27_DFFPOSX1_17 ( );
FILL FILL_0_DFFPOSX1_24 ( );
FILL FILL_1_DFFPOSX1_24 ( );
FILL FILL_2_DFFPOSX1_24 ( );
FILL FILL_3_DFFPOSX1_24 ( );
FILL FILL_4_DFFPOSX1_24 ( );
FILL FILL_5_DFFPOSX1_24 ( );
FILL FILL_6_DFFPOSX1_24 ( );
FILL FILL_7_DFFPOSX1_24 ( );
FILL FILL_8_DFFPOSX1_24 ( );
FILL FILL_9_DFFPOSX1_24 ( );
FILL FILL_10_DFFPOSX1_24 ( );
FILL FILL_11_DFFPOSX1_24 ( );
FILL FILL_12_DFFPOSX1_24 ( );
FILL FILL_13_DFFPOSX1_24 ( );
FILL FILL_14_DFFPOSX1_24 ( );
FILL FILL_15_DFFPOSX1_24 ( );
FILL FILL_16_DFFPOSX1_24 ( );
FILL FILL_17_DFFPOSX1_24 ( );
FILL FILL_18_DFFPOSX1_24 ( );
FILL FILL_19_DFFPOSX1_24 ( );
FILL FILL_20_DFFPOSX1_24 ( );
FILL FILL_21_DFFPOSX1_24 ( );
FILL FILL_22_DFFPOSX1_24 ( );
FILL FILL_23_DFFPOSX1_24 ( );
FILL FILL_24_DFFPOSX1_24 ( );
FILL FILL_25_DFFPOSX1_24 ( );
FILL FILL_26_DFFPOSX1_24 ( );
FILL FILL_27_DFFPOSX1_24 ( );
FILL FILL_0_NOR2X1_75 ( );
FILL FILL_1_NOR2X1_75 ( );
FILL FILL_2_NOR2X1_75 ( );
FILL FILL_3_NOR2X1_75 ( );
FILL FILL_4_NOR2X1_75 ( );
FILL FILL_5_NOR2X1_75 ( );
FILL FILL_6_NOR2X1_75 ( );
FILL FILL_0_INVX1_130 ( );
FILL FILL_1_INVX1_130 ( );
FILL FILL_2_INVX1_130 ( );
FILL FILL_3_INVX1_130 ( );
FILL FILL_4_INVX1_130 ( );
FILL FILL_0_AND2X2_28 ( );
FILL FILL_1_AND2X2_28 ( );
FILL FILL_2_AND2X2_28 ( );
FILL FILL_3_AND2X2_28 ( );
FILL FILL_4_AND2X2_28 ( );
FILL FILL_5_AND2X2_28 ( );
FILL FILL_6_AND2X2_28 ( );
FILL FILL_7_AND2X2_28 ( );
FILL FILL_8_AND2X2_28 ( );
FILL FILL_9_AND2X2_28 ( );
FILL FILL_0_BUFX2_8 ( );
FILL FILL_1_BUFX2_8 ( );
FILL FILL_2_BUFX2_8 ( );
FILL FILL_3_BUFX2_8 ( );
FILL FILL_4_BUFX2_8 ( );
FILL FILL_5_BUFX2_8 ( );
FILL FILL_6_BUFX2_8 ( );
FILL FILL_0_OAI21X1_91 ( );
FILL FILL_1_OAI21X1_91 ( );
FILL FILL_2_OAI21X1_91 ( );
FILL FILL_3_OAI21X1_91 ( );
FILL FILL_4_OAI21X1_91 ( );
FILL FILL_5_OAI21X1_91 ( );
FILL FILL_6_OAI21X1_91 ( );
FILL FILL_7_OAI21X1_91 ( );
FILL FILL_8_OAI21X1_91 ( );
FILL FILL_0_DFFSR_51 ( );
FILL FILL_1_DFFSR_51 ( );
FILL FILL_2_DFFSR_51 ( );
FILL FILL_3_DFFSR_51 ( );
FILL FILL_4_DFFSR_51 ( );
FILL FILL_5_DFFSR_51 ( );
FILL FILL_6_DFFSR_51 ( );
FILL FILL_7_DFFSR_51 ( );
FILL FILL_8_DFFSR_51 ( );
FILL FILL_9_DFFSR_51 ( );
FILL FILL_10_DFFSR_51 ( );
FILL FILL_11_DFFSR_51 ( );
FILL FILL_12_DFFSR_51 ( );
FILL FILL_13_DFFSR_51 ( );
FILL FILL_14_DFFSR_51 ( );
FILL FILL_15_DFFSR_51 ( );
FILL FILL_16_DFFSR_51 ( );
FILL FILL_17_DFFSR_51 ( );
FILL FILL_18_DFFSR_51 ( );
FILL FILL_19_DFFSR_51 ( );
FILL FILL_20_DFFSR_51 ( );
FILL FILL_21_DFFSR_51 ( );
FILL FILL_22_DFFSR_51 ( );
FILL FILL_23_DFFSR_51 ( );
FILL FILL_24_DFFSR_51 ( );
FILL FILL_25_DFFSR_51 ( );
FILL FILL_26_DFFSR_51 ( );
FILL FILL_27_DFFSR_51 ( );
FILL FILL_28_DFFSR_51 ( );
FILL FILL_29_DFFSR_51 ( );
FILL FILL_30_DFFSR_51 ( );
FILL FILL_31_DFFSR_51 ( );
FILL FILL_32_DFFSR_51 ( );
FILL FILL_33_DFFSR_51 ( );
FILL FILL_34_DFFSR_51 ( );
FILL FILL_35_DFFSR_51 ( );
FILL FILL_36_DFFSR_51 ( );
FILL FILL_37_DFFSR_51 ( );
FILL FILL_38_DFFSR_51 ( );
FILL FILL_39_DFFSR_51 ( );
FILL FILL_40_DFFSR_51 ( );
FILL FILL_41_DFFSR_51 ( );
FILL FILL_42_DFFSR_51 ( );
FILL FILL_43_DFFSR_51 ( );
FILL FILL_44_DFFSR_51 ( );
FILL FILL_45_DFFSR_51 ( );
FILL FILL_46_DFFSR_51 ( );
FILL FILL_47_DFFSR_51 ( );
FILL FILL_48_DFFSR_51 ( );
FILL FILL_49_DFFSR_51 ( );
FILL FILL_50_DFFSR_51 ( );
FILL FILL_51_DFFSR_51 ( );
FILL FILL_0_CLKBUF1_11 ( );
FILL FILL_1_CLKBUF1_11 ( );
FILL FILL_2_CLKBUF1_11 ( );
FILL FILL_3_CLKBUF1_11 ( );
FILL FILL_4_CLKBUF1_11 ( );
FILL FILL_5_CLKBUF1_11 ( );
FILL FILL_6_CLKBUF1_11 ( );
FILL FILL_7_CLKBUF1_11 ( );
FILL FILL_8_CLKBUF1_11 ( );
FILL FILL_9_CLKBUF1_11 ( );
FILL FILL_10_CLKBUF1_11 ( );
FILL FILL_11_CLKBUF1_11 ( );
FILL FILL_12_CLKBUF1_11 ( );
FILL FILL_13_CLKBUF1_11 ( );
FILL FILL_14_CLKBUF1_11 ( );
FILL FILL_15_CLKBUF1_11 ( );
FILL FILL_16_CLKBUF1_11 ( );
FILL FILL_17_CLKBUF1_11 ( );
FILL FILL_18_CLKBUF1_11 ( );
FILL FILL_19_CLKBUF1_11 ( );
FILL FILL_20_CLKBUF1_11 ( );
FILL FILL_0_NOR2X1_61 ( );
FILL FILL_1_NOR2X1_61 ( );
FILL FILL_2_NOR2X1_61 ( );
FILL FILL_3_NOR2X1_61 ( );
FILL FILL_4_NOR2X1_61 ( );
FILL FILL_5_NOR2X1_61 ( );
FILL FILL_6_NOR2X1_61 ( );
FILL FILL_0_INVX1_127 ( );
FILL FILL_1_INVX1_127 ( );
FILL FILL_2_INVX1_127 ( );
FILL FILL_3_INVX1_127 ( );
FILL FILL_4_INVX1_127 ( );
FILL FILL_0_NAND3X1_133 ( );
FILL FILL_1_NAND3X1_133 ( );
FILL FILL_2_NAND3X1_133 ( );
FILL FILL_3_NAND3X1_133 ( );
FILL FILL_4_NAND3X1_133 ( );
FILL FILL_5_NAND3X1_133 ( );
FILL FILL_6_NAND3X1_133 ( );
FILL FILL_7_NAND3X1_133 ( );
FILL FILL_8_NAND3X1_133 ( );
FILL FILL_0_DFFSR_174 ( );
FILL FILL_1_DFFSR_174 ( );
FILL FILL_2_DFFSR_174 ( );
FILL FILL_3_DFFSR_174 ( );
FILL FILL_4_DFFSR_174 ( );
FILL FILL_5_DFFSR_174 ( );
FILL FILL_6_DFFSR_174 ( );
FILL FILL_7_DFFSR_174 ( );
FILL FILL_8_DFFSR_174 ( );
FILL FILL_9_DFFSR_174 ( );
FILL FILL_10_DFFSR_174 ( );
FILL FILL_11_DFFSR_174 ( );
FILL FILL_12_DFFSR_174 ( );
FILL FILL_13_DFFSR_174 ( );
FILL FILL_14_DFFSR_174 ( );
FILL FILL_15_DFFSR_174 ( );
FILL FILL_16_DFFSR_174 ( );
FILL FILL_17_DFFSR_174 ( );
FILL FILL_18_DFFSR_174 ( );
FILL FILL_19_DFFSR_174 ( );
FILL FILL_20_DFFSR_174 ( );
FILL FILL_21_DFFSR_174 ( );
FILL FILL_22_DFFSR_174 ( );
FILL FILL_23_DFFSR_174 ( );
FILL FILL_24_DFFSR_174 ( );
FILL FILL_25_DFFSR_174 ( );
FILL FILL_26_DFFSR_174 ( );
FILL FILL_27_DFFSR_174 ( );
FILL FILL_28_DFFSR_174 ( );
FILL FILL_29_DFFSR_174 ( );
FILL FILL_30_DFFSR_174 ( );
FILL FILL_31_DFFSR_174 ( );
FILL FILL_32_DFFSR_174 ( );
FILL FILL_33_DFFSR_174 ( );
FILL FILL_34_DFFSR_174 ( );
FILL FILL_35_DFFSR_174 ( );
FILL FILL_36_DFFSR_174 ( );
FILL FILL_37_DFFSR_174 ( );
FILL FILL_38_DFFSR_174 ( );
FILL FILL_39_DFFSR_174 ( );
FILL FILL_40_DFFSR_174 ( );
FILL FILL_41_DFFSR_174 ( );
FILL FILL_42_DFFSR_174 ( );
FILL FILL_43_DFFSR_174 ( );
FILL FILL_44_DFFSR_174 ( );
FILL FILL_45_DFFSR_174 ( );
FILL FILL_46_DFFSR_174 ( );
FILL FILL_47_DFFSR_174 ( );
FILL FILL_48_DFFSR_174 ( );
FILL FILL_49_DFFSR_174 ( );
FILL FILL_50_DFFSR_174 ( );
FILL FILL_0_AND2X2_24 ( );
FILL FILL_1_AND2X2_24 ( );
FILL FILL_2_AND2X2_24 ( );
FILL FILL_3_AND2X2_24 ( );
FILL FILL_4_AND2X2_24 ( );
FILL FILL_5_AND2X2_24 ( );
FILL FILL_6_AND2X2_24 ( );
FILL FILL_7_AND2X2_24 ( );
FILL FILL_8_AND2X2_24 ( );
FILL FILL_0_OAI22X1_42 ( );
FILL FILL_1_OAI22X1_42 ( );
FILL FILL_2_OAI22X1_42 ( );
FILL FILL_3_OAI22X1_42 ( );
FILL FILL_4_OAI22X1_42 ( );
FILL FILL_5_OAI22X1_42 ( );
FILL FILL_6_OAI22X1_42 ( );
FILL FILL_7_OAI22X1_42 ( );
FILL FILL_8_OAI22X1_42 ( );
FILL FILL_9_OAI22X1_42 ( );
FILL FILL_10_OAI22X1_42 ( );
FILL FILL_11_OAI22X1_42 ( );
FILL FILL_0_BUFX2_29 ( );
FILL FILL_1_BUFX2_29 ( );
FILL FILL_2_BUFX2_29 ( );
FILL FILL_3_BUFX2_29 ( );
FILL FILL_4_BUFX2_29 ( );
FILL FILL_5_BUFX2_29 ( );
FILL FILL_6_BUFX2_29 ( );
FILL FILL_0_BUFX2_32 ( );
FILL FILL_1_BUFX2_32 ( );
FILL FILL_2_BUFX2_32 ( );
FILL FILL_3_BUFX2_32 ( );
FILL FILL_4_BUFX2_32 ( );
FILL FILL_5_BUFX2_32 ( );
FILL FILL_6_BUFX2_32 ( );
FILL FILL_0_BUFX2_26 ( );
FILL FILL_1_BUFX2_26 ( );
FILL FILL_2_BUFX2_26 ( );
FILL FILL_3_BUFX2_26 ( );
FILL FILL_4_BUFX2_26 ( );
FILL FILL_5_BUFX2_26 ( );
FILL FILL_6_BUFX2_26 ( );
FILL FILL_0_CLKBUF1_20 ( );
FILL FILL_1_CLKBUF1_20 ( );
FILL FILL_2_CLKBUF1_20 ( );
FILL FILL_3_CLKBUF1_20 ( );
FILL FILL_4_CLKBUF1_20 ( );
FILL FILL_5_CLKBUF1_20 ( );
FILL FILL_6_CLKBUF1_20 ( );
FILL FILL_7_CLKBUF1_20 ( );
FILL FILL_8_CLKBUF1_20 ( );
FILL FILL_9_CLKBUF1_20 ( );
FILL FILL_10_CLKBUF1_20 ( );
FILL FILL_11_CLKBUF1_20 ( );
FILL FILL_12_CLKBUF1_20 ( );
FILL FILL_13_CLKBUF1_20 ( );
FILL FILL_14_CLKBUF1_20 ( );
FILL FILL_15_CLKBUF1_20 ( );
FILL FILL_16_CLKBUF1_20 ( );
FILL FILL_17_CLKBUF1_20 ( );
FILL FILL_18_CLKBUF1_20 ( );
FILL FILL_19_CLKBUF1_20 ( );
FILL FILL_20_CLKBUF1_20 ( );
FILL FILL_21_CLKBUF1_20 ( );
FILL FILL_0_BUFX2_94 ( );
FILL FILL_1_BUFX2_94 ( );
FILL FILL_2_BUFX2_94 ( );
FILL FILL_3_BUFX2_94 ( );
FILL FILL_4_BUFX2_94 ( );
FILL FILL_5_BUFX2_94 ( );
FILL FILL_6_BUFX2_94 ( );
FILL FILL_0_NAND3X1_120 ( );
FILL FILL_1_NAND3X1_120 ( );
FILL FILL_2_NAND3X1_120 ( );
FILL FILL_3_NAND3X1_120 ( );
FILL FILL_4_NAND3X1_120 ( );
FILL FILL_5_NAND3X1_120 ( );
FILL FILL_6_NAND3X1_120 ( );
FILL FILL_7_NAND3X1_120 ( );
FILL FILL_8_NAND3X1_120 ( );
FILL FILL_0_NOR2X1_54 ( );
FILL FILL_1_NOR2X1_54 ( );
FILL FILL_2_NOR2X1_54 ( );
FILL FILL_3_NOR2X1_54 ( );
FILL FILL_4_NOR2X1_54 ( );
FILL FILL_5_NOR2X1_54 ( );
FILL FILL_6_NOR2X1_54 ( );
FILL FILL_0_DFFSR_189 ( );
FILL FILL_1_DFFSR_189 ( );
FILL FILL_2_DFFSR_189 ( );
FILL FILL_3_DFFSR_189 ( );
FILL FILL_4_DFFSR_189 ( );
FILL FILL_5_DFFSR_189 ( );
FILL FILL_6_DFFSR_189 ( );
FILL FILL_7_DFFSR_189 ( );
FILL FILL_8_DFFSR_189 ( );
FILL FILL_9_DFFSR_189 ( );
FILL FILL_10_DFFSR_189 ( );
FILL FILL_11_DFFSR_189 ( );
FILL FILL_12_DFFSR_189 ( );
FILL FILL_13_DFFSR_189 ( );
FILL FILL_14_DFFSR_189 ( );
FILL FILL_15_DFFSR_189 ( );
FILL FILL_16_DFFSR_189 ( );
FILL FILL_17_DFFSR_189 ( );
FILL FILL_18_DFFSR_189 ( );
FILL FILL_19_DFFSR_189 ( );
FILL FILL_20_DFFSR_189 ( );
FILL FILL_21_DFFSR_189 ( );
FILL FILL_22_DFFSR_189 ( );
FILL FILL_23_DFFSR_189 ( );
FILL FILL_24_DFFSR_189 ( );
FILL FILL_25_DFFSR_189 ( );
FILL FILL_26_DFFSR_189 ( );
FILL FILL_27_DFFSR_189 ( );
FILL FILL_28_DFFSR_189 ( );
FILL FILL_29_DFFSR_189 ( );
FILL FILL_30_DFFSR_189 ( );
FILL FILL_31_DFFSR_189 ( );
FILL FILL_32_DFFSR_189 ( );
FILL FILL_33_DFFSR_189 ( );
FILL FILL_34_DFFSR_189 ( );
FILL FILL_35_DFFSR_189 ( );
FILL FILL_36_DFFSR_189 ( );
FILL FILL_37_DFFSR_189 ( );
FILL FILL_38_DFFSR_189 ( );
FILL FILL_39_DFFSR_189 ( );
FILL FILL_40_DFFSR_189 ( );
FILL FILL_41_DFFSR_189 ( );
FILL FILL_42_DFFSR_189 ( );
FILL FILL_43_DFFSR_189 ( );
FILL FILL_44_DFFSR_189 ( );
FILL FILL_45_DFFSR_189 ( );
FILL FILL_46_DFFSR_189 ( );
FILL FILL_47_DFFSR_189 ( );
FILL FILL_48_DFFSR_189 ( );
FILL FILL_49_DFFSR_189 ( );
FILL FILL_50_DFFSR_189 ( );
FILL FILL_0_NAND2X1_102 ( );
FILL FILL_1_NAND2X1_102 ( );
FILL FILL_2_NAND2X1_102 ( );
FILL FILL_3_NAND2X1_102 ( );
FILL FILL_4_NAND2X1_102 ( );
FILL FILL_5_NAND2X1_102 ( );
FILL FILL_6_NAND2X1_102 ( );
FILL FILL_0_OAI21X1_60 ( );
FILL FILL_1_OAI21X1_60 ( );
FILL FILL_2_OAI21X1_60 ( );
FILL FILL_3_OAI21X1_60 ( );
FILL FILL_4_OAI21X1_60 ( );
FILL FILL_5_OAI21X1_60 ( );
FILL FILL_6_OAI21X1_60 ( );
FILL FILL_7_OAI21X1_60 ( );
FILL FILL_8_OAI21X1_60 ( );
FILL FILL_0_AOI21X1_27 ( );
FILL FILL_1_AOI21X1_27 ( );
FILL FILL_2_AOI21X1_27 ( );
FILL FILL_3_AOI21X1_27 ( );
FILL FILL_4_AOI21X1_27 ( );
FILL FILL_5_AOI21X1_27 ( );
FILL FILL_6_AOI21X1_27 ( );
FILL FILL_7_AOI21X1_27 ( );
FILL FILL_8_AOI21X1_27 ( );
FILL FILL_0_INVX1_133 ( );
FILL FILL_1_INVX1_133 ( );
FILL FILL_2_INVX1_133 ( );
FILL FILL_3_INVX1_133 ( );
FILL FILL_4_INVX1_133 ( );
FILL FILL_0_INVX1_151 ( );
FILL FILL_1_INVX1_151 ( );
FILL FILL_2_INVX1_151 ( );
FILL FILL_3_INVX1_151 ( );
FILL FILL_0_NAND3X1_160 ( );
FILL FILL_1_NAND3X1_160 ( );
FILL FILL_2_NAND3X1_160 ( );
FILL FILL_3_NAND3X1_160 ( );
FILL FILL_4_NAND3X1_160 ( );
FILL FILL_5_NAND3X1_160 ( );
FILL FILL_6_NAND3X1_160 ( );
FILL FILL_7_NAND3X1_160 ( );
FILL FILL_8_NAND3X1_160 ( );
FILL FILL_0_AOI21X1_11 ( );
FILL FILL_1_AOI21X1_11 ( );
FILL FILL_2_AOI21X1_11 ( );
FILL FILL_3_AOI21X1_11 ( );
FILL FILL_4_AOI21X1_11 ( );
FILL FILL_5_AOI21X1_11 ( );
FILL FILL_6_AOI21X1_11 ( );
FILL FILL_7_AOI21X1_11 ( );
FILL FILL_8_AOI21X1_11 ( );
FILL FILL_9_AOI21X1_11 ( );
FILL FILL_0_INVX1_145 ( );
FILL FILL_1_INVX1_145 ( );
FILL FILL_2_INVX1_145 ( );
FILL FILL_3_INVX1_145 ( );
FILL FILL_4_INVX1_145 ( );
FILL FILL_0_NAND3X1_147 ( );
FILL FILL_1_NAND3X1_147 ( );
FILL FILL_2_NAND3X1_147 ( );
FILL FILL_3_NAND3X1_147 ( );
FILL FILL_4_NAND3X1_147 ( );
FILL FILL_5_NAND3X1_147 ( );
FILL FILL_6_NAND3X1_147 ( );
FILL FILL_7_NAND3X1_147 ( );
FILL FILL_8_NAND3X1_147 ( );
FILL FILL_0_AOI22X1_19 ( );
FILL FILL_1_AOI22X1_19 ( );
FILL FILL_2_AOI22X1_19 ( );
FILL FILL_3_AOI22X1_19 ( );
FILL FILL_4_AOI22X1_19 ( );
FILL FILL_5_AOI22X1_19 ( );
FILL FILL_6_AOI22X1_19 ( );
FILL FILL_7_AOI22X1_19 ( );
FILL FILL_8_AOI22X1_19 ( );
FILL FILL_9_AOI22X1_19 ( );
FILL FILL_10_AOI22X1_19 ( );
FILL FILL_11_AOI22X1_19 ( );
FILL FILL_0_NAND2X1_127 ( );
FILL FILL_1_NAND2X1_127 ( );
FILL FILL_2_NAND2X1_127 ( );
FILL FILL_3_NAND2X1_127 ( );
FILL FILL_4_NAND2X1_127 ( );
FILL FILL_5_NAND2X1_127 ( );
FILL FILL_6_NAND2X1_127 ( );
FILL FILL_0_DFFSR_268 ( );
FILL FILL_1_DFFSR_268 ( );
FILL FILL_2_DFFSR_268 ( );
FILL FILL_3_DFFSR_268 ( );
FILL FILL_4_DFFSR_268 ( );
FILL FILL_5_DFFSR_268 ( );
FILL FILL_6_DFFSR_268 ( );
FILL FILL_7_DFFSR_268 ( );
FILL FILL_8_DFFSR_268 ( );
FILL FILL_9_DFFSR_268 ( );
FILL FILL_10_DFFSR_268 ( );
FILL FILL_11_DFFSR_268 ( );
FILL FILL_12_DFFSR_268 ( );
FILL FILL_13_DFFSR_268 ( );
FILL FILL_14_DFFSR_268 ( );
FILL FILL_15_DFFSR_268 ( );
FILL FILL_16_DFFSR_268 ( );
FILL FILL_17_DFFSR_268 ( );
FILL FILL_18_DFFSR_268 ( );
FILL FILL_19_DFFSR_268 ( );
FILL FILL_20_DFFSR_268 ( );
FILL FILL_21_DFFSR_268 ( );
FILL FILL_22_DFFSR_268 ( );
FILL FILL_23_DFFSR_268 ( );
FILL FILL_24_DFFSR_268 ( );
FILL FILL_25_DFFSR_268 ( );
FILL FILL_26_DFFSR_268 ( );
FILL FILL_27_DFFSR_268 ( );
FILL FILL_28_DFFSR_268 ( );
FILL FILL_29_DFFSR_268 ( );
FILL FILL_30_DFFSR_268 ( );
FILL FILL_31_DFFSR_268 ( );
FILL FILL_32_DFFSR_268 ( );
FILL FILL_33_DFFSR_268 ( );
FILL FILL_34_DFFSR_268 ( );
FILL FILL_35_DFFSR_268 ( );
FILL FILL_36_DFFSR_268 ( );
FILL FILL_37_DFFSR_268 ( );
FILL FILL_38_DFFSR_268 ( );
FILL FILL_39_DFFSR_268 ( );
FILL FILL_40_DFFSR_268 ( );
FILL FILL_41_DFFSR_268 ( );
FILL FILL_42_DFFSR_268 ( );
FILL FILL_43_DFFSR_268 ( );
FILL FILL_44_DFFSR_268 ( );
FILL FILL_45_DFFSR_268 ( );
FILL FILL_46_DFFSR_268 ( );
FILL FILL_47_DFFSR_268 ( );
FILL FILL_48_DFFSR_268 ( );
FILL FILL_49_DFFSR_268 ( );
FILL FILL_50_DFFSR_268 ( );
FILL FILL_51_DFFSR_268 ( );
FILL FILL_0_AOI21X1_59 ( );
FILL FILL_1_AOI21X1_59 ( );
FILL FILL_2_AOI21X1_59 ( );
FILL FILL_3_AOI21X1_59 ( );
FILL FILL_4_AOI21X1_59 ( );
FILL FILL_5_AOI21X1_59 ( );
FILL FILL_6_AOI21X1_59 ( );
FILL FILL_7_AOI21X1_59 ( );
FILL FILL_8_AOI21X1_59 ( );
FILL FILL_9_AOI21X1_59 ( );
FILL FILL_0_DFFPOSX1_38 ( );
FILL FILL_1_DFFPOSX1_38 ( );
FILL FILL_2_DFFPOSX1_38 ( );
FILL FILL_3_DFFPOSX1_38 ( );
FILL FILL_4_DFFPOSX1_38 ( );
FILL FILL_5_DFFPOSX1_38 ( );
FILL FILL_6_DFFPOSX1_38 ( );
FILL FILL_7_DFFPOSX1_38 ( );
FILL FILL_8_DFFPOSX1_38 ( );
FILL FILL_9_DFFPOSX1_38 ( );
FILL FILL_10_DFFPOSX1_38 ( );
FILL FILL_11_DFFPOSX1_38 ( );
FILL FILL_12_DFFPOSX1_38 ( );
FILL FILL_13_DFFPOSX1_38 ( );
FILL FILL_14_DFFPOSX1_38 ( );
FILL FILL_15_DFFPOSX1_38 ( );
FILL FILL_16_DFFPOSX1_38 ( );
FILL FILL_17_DFFPOSX1_38 ( );
FILL FILL_18_DFFPOSX1_38 ( );
FILL FILL_19_DFFPOSX1_38 ( );
FILL FILL_20_DFFPOSX1_38 ( );
FILL FILL_21_DFFPOSX1_38 ( );
FILL FILL_22_DFFPOSX1_38 ( );
FILL FILL_23_DFFPOSX1_38 ( );
FILL FILL_24_DFFPOSX1_38 ( );
FILL FILL_25_DFFPOSX1_38 ( );
FILL FILL_26_DFFPOSX1_38 ( );
FILL FILL_27_DFFPOSX1_38 ( );
FILL FILL_0_DFFSR_263 ( );
FILL FILL_1_DFFSR_263 ( );
FILL FILL_2_DFFSR_263 ( );
FILL FILL_3_DFFSR_263 ( );
FILL FILL_4_DFFSR_263 ( );
FILL FILL_5_DFFSR_263 ( );
FILL FILL_6_DFFSR_263 ( );
FILL FILL_7_DFFSR_263 ( );
FILL FILL_8_DFFSR_263 ( );
FILL FILL_9_DFFSR_263 ( );
FILL FILL_10_DFFSR_263 ( );
FILL FILL_11_DFFSR_263 ( );
FILL FILL_12_DFFSR_263 ( );
FILL FILL_13_DFFSR_263 ( );
FILL FILL_14_DFFSR_263 ( );
FILL FILL_15_DFFSR_263 ( );
FILL FILL_16_DFFSR_263 ( );
FILL FILL_17_DFFSR_263 ( );
FILL FILL_18_DFFSR_263 ( );
FILL FILL_19_DFFSR_263 ( );
FILL FILL_20_DFFSR_263 ( );
FILL FILL_21_DFFSR_263 ( );
FILL FILL_22_DFFSR_263 ( );
FILL FILL_23_DFFSR_263 ( );
FILL FILL_24_DFFSR_263 ( );
FILL FILL_25_DFFSR_263 ( );
FILL FILL_26_DFFSR_263 ( );
FILL FILL_27_DFFSR_263 ( );
FILL FILL_28_DFFSR_263 ( );
FILL FILL_29_DFFSR_263 ( );
FILL FILL_30_DFFSR_263 ( );
FILL FILL_31_DFFSR_263 ( );
FILL FILL_32_DFFSR_263 ( );
FILL FILL_33_DFFSR_263 ( );
FILL FILL_34_DFFSR_263 ( );
FILL FILL_35_DFFSR_263 ( );
FILL FILL_36_DFFSR_263 ( );
FILL FILL_37_DFFSR_263 ( );
FILL FILL_38_DFFSR_263 ( );
FILL FILL_39_DFFSR_263 ( );
FILL FILL_40_DFFSR_263 ( );
FILL FILL_41_DFFSR_263 ( );
FILL FILL_42_DFFSR_263 ( );
FILL FILL_43_DFFSR_263 ( );
FILL FILL_44_DFFSR_263 ( );
FILL FILL_45_DFFSR_263 ( );
FILL FILL_46_DFFSR_263 ( );
FILL FILL_47_DFFSR_263 ( );
FILL FILL_48_DFFSR_263 ( );
FILL FILL_49_DFFSR_263 ( );
FILL FILL_50_DFFSR_263 ( );
FILL FILL_0_CLKBUF1_18 ( );
FILL FILL_1_CLKBUF1_18 ( );
FILL FILL_2_CLKBUF1_18 ( );
FILL FILL_3_CLKBUF1_18 ( );
FILL FILL_4_CLKBUF1_18 ( );
FILL FILL_5_CLKBUF1_18 ( );
FILL FILL_6_CLKBUF1_18 ( );
FILL FILL_7_CLKBUF1_18 ( );
FILL FILL_8_CLKBUF1_18 ( );
FILL FILL_9_CLKBUF1_18 ( );
FILL FILL_10_CLKBUF1_18 ( );
FILL FILL_11_CLKBUF1_18 ( );
FILL FILL_12_CLKBUF1_18 ( );
FILL FILL_13_CLKBUF1_18 ( );
FILL FILL_14_CLKBUF1_18 ( );
FILL FILL_15_CLKBUF1_18 ( );
FILL FILL_16_CLKBUF1_18 ( );
FILL FILL_17_CLKBUF1_18 ( );
FILL FILL_18_CLKBUF1_18 ( );
FILL FILL_19_CLKBUF1_18 ( );
FILL FILL_20_CLKBUF1_18 ( );
FILL FILL_0_DFFSR_73 ( );
FILL FILL_1_DFFSR_73 ( );
FILL FILL_2_DFFSR_73 ( );
FILL FILL_3_DFFSR_73 ( );
FILL FILL_4_DFFSR_73 ( );
FILL FILL_5_DFFSR_73 ( );
FILL FILL_6_DFFSR_73 ( );
FILL FILL_7_DFFSR_73 ( );
FILL FILL_8_DFFSR_73 ( );
FILL FILL_9_DFFSR_73 ( );
FILL FILL_10_DFFSR_73 ( );
FILL FILL_11_DFFSR_73 ( );
FILL FILL_12_DFFSR_73 ( );
FILL FILL_13_DFFSR_73 ( );
FILL FILL_14_DFFSR_73 ( );
FILL FILL_15_DFFSR_73 ( );
FILL FILL_16_DFFSR_73 ( );
FILL FILL_17_DFFSR_73 ( );
FILL FILL_18_DFFSR_73 ( );
FILL FILL_19_DFFSR_73 ( );
FILL FILL_20_DFFSR_73 ( );
FILL FILL_21_DFFSR_73 ( );
FILL FILL_22_DFFSR_73 ( );
FILL FILL_23_DFFSR_73 ( );
FILL FILL_24_DFFSR_73 ( );
FILL FILL_25_DFFSR_73 ( );
FILL FILL_26_DFFSR_73 ( );
FILL FILL_27_DFFSR_73 ( );
FILL FILL_28_DFFSR_73 ( );
FILL FILL_29_DFFSR_73 ( );
FILL FILL_30_DFFSR_73 ( );
FILL FILL_31_DFFSR_73 ( );
FILL FILL_32_DFFSR_73 ( );
FILL FILL_33_DFFSR_73 ( );
FILL FILL_34_DFFSR_73 ( );
FILL FILL_35_DFFSR_73 ( );
FILL FILL_36_DFFSR_73 ( );
FILL FILL_37_DFFSR_73 ( );
FILL FILL_38_DFFSR_73 ( );
FILL FILL_39_DFFSR_73 ( );
FILL FILL_40_DFFSR_73 ( );
FILL FILL_41_DFFSR_73 ( );
FILL FILL_42_DFFSR_73 ( );
FILL FILL_43_DFFSR_73 ( );
FILL FILL_44_DFFSR_73 ( );
FILL FILL_45_DFFSR_73 ( );
FILL FILL_46_DFFSR_73 ( );
FILL FILL_47_DFFSR_73 ( );
FILL FILL_48_DFFSR_73 ( );
FILL FILL_49_DFFSR_73 ( );
FILL FILL_50_DFFSR_73 ( );
FILL FILL_0_INVX1_89 ( );
FILL FILL_1_INVX1_89 ( );
FILL FILL_2_INVX1_89 ( );
FILL FILL_3_INVX1_89 ( );
FILL FILL_0_OAI21X1_12 ( );
FILL FILL_1_OAI21X1_12 ( );
FILL FILL_2_OAI21X1_12 ( );
FILL FILL_3_OAI21X1_12 ( );
FILL FILL_4_OAI21X1_12 ( );
FILL FILL_5_OAI21X1_12 ( );
FILL FILL_6_OAI21X1_12 ( );
FILL FILL_7_OAI21X1_12 ( );
FILL FILL_8_OAI21X1_12 ( );
FILL FILL_9_OAI21X1_12 ( );
FILL FILL_0_NOR2X1_36 ( );
FILL FILL_1_NOR2X1_36 ( );
FILL FILL_2_NOR2X1_36 ( );
FILL FILL_3_NOR2X1_36 ( );
FILL FILL_4_NOR2X1_36 ( );
FILL FILL_5_NOR2X1_36 ( );
FILL FILL_6_NOR2X1_36 ( );
FILL FILL_0_INVX1_81 ( );
FILL FILL_1_INVX1_81 ( );
FILL FILL_2_INVX1_81 ( );
FILL FILL_3_INVX1_81 ( );
FILL FILL_0_OAI22X1_33 ( );
FILL FILL_1_OAI22X1_33 ( );
FILL FILL_2_OAI22X1_33 ( );
FILL FILL_3_OAI22X1_33 ( );
FILL FILL_4_OAI22X1_33 ( );
FILL FILL_5_OAI22X1_33 ( );
FILL FILL_6_OAI22X1_33 ( );
FILL FILL_7_OAI22X1_33 ( );
FILL FILL_8_OAI22X1_33 ( );
FILL FILL_9_OAI22X1_33 ( );
FILL FILL_10_OAI22X1_33 ( );
FILL FILL_11_OAI22X1_33 ( );
FILL FILL_0_INVX1_101 ( );
FILL FILL_1_INVX1_101 ( );
FILL FILL_2_INVX1_101 ( );
FILL FILL_3_INVX1_101 ( );
FILL FILL_4_INVX1_101 ( );
FILL FILL_0_DFFSR_179 ( );
FILL FILL_1_DFFSR_179 ( );
FILL FILL_2_DFFSR_179 ( );
FILL FILL_3_DFFSR_179 ( );
FILL FILL_4_DFFSR_179 ( );
FILL FILL_5_DFFSR_179 ( );
FILL FILL_6_DFFSR_179 ( );
FILL FILL_7_DFFSR_179 ( );
FILL FILL_8_DFFSR_179 ( );
FILL FILL_9_DFFSR_179 ( );
FILL FILL_10_DFFSR_179 ( );
FILL FILL_11_DFFSR_179 ( );
FILL FILL_12_DFFSR_179 ( );
FILL FILL_13_DFFSR_179 ( );
FILL FILL_14_DFFSR_179 ( );
FILL FILL_15_DFFSR_179 ( );
FILL FILL_16_DFFSR_179 ( );
FILL FILL_17_DFFSR_179 ( );
FILL FILL_18_DFFSR_179 ( );
FILL FILL_19_DFFSR_179 ( );
FILL FILL_20_DFFSR_179 ( );
FILL FILL_21_DFFSR_179 ( );
FILL FILL_22_DFFSR_179 ( );
FILL FILL_23_DFFSR_179 ( );
FILL FILL_24_DFFSR_179 ( );
FILL FILL_25_DFFSR_179 ( );
FILL FILL_26_DFFSR_179 ( );
FILL FILL_27_DFFSR_179 ( );
FILL FILL_28_DFFSR_179 ( );
FILL FILL_29_DFFSR_179 ( );
FILL FILL_30_DFFSR_179 ( );
FILL FILL_31_DFFSR_179 ( );
FILL FILL_32_DFFSR_179 ( );
FILL FILL_33_DFFSR_179 ( );
FILL FILL_34_DFFSR_179 ( );
FILL FILL_35_DFFSR_179 ( );
FILL FILL_36_DFFSR_179 ( );
FILL FILL_37_DFFSR_179 ( );
FILL FILL_38_DFFSR_179 ( );
FILL FILL_39_DFFSR_179 ( );
FILL FILL_40_DFFSR_179 ( );
FILL FILL_41_DFFSR_179 ( );
FILL FILL_42_DFFSR_179 ( );
FILL FILL_43_DFFSR_179 ( );
FILL FILL_44_DFFSR_179 ( );
FILL FILL_45_DFFSR_179 ( );
FILL FILL_46_DFFSR_179 ( );
FILL FILL_47_DFFSR_179 ( );
FILL FILL_48_DFFSR_179 ( );
FILL FILL_49_DFFSR_179 ( );
FILL FILL_50_DFFSR_179 ( );
FILL FILL_51_DFFSR_179 ( );
FILL FILL_0_NAND3X1_99 ( );
FILL FILL_1_NAND3X1_99 ( );
FILL FILL_2_NAND3X1_99 ( );
FILL FILL_3_NAND3X1_99 ( );
FILL FILL_4_NAND3X1_99 ( );
FILL FILL_5_NAND3X1_99 ( );
FILL FILL_6_NAND3X1_99 ( );
FILL FILL_7_NAND3X1_99 ( );
FILL FILL_8_NAND3X1_99 ( );
FILL FILL_0_BUFX2_30 ( );
FILL FILL_1_BUFX2_30 ( );
FILL FILL_2_BUFX2_30 ( );
FILL FILL_3_BUFX2_30 ( );
FILL FILL_4_BUFX2_30 ( );
FILL FILL_5_BUFX2_30 ( );
FILL FILL_6_BUFX2_30 ( );
FILL FILL_0_DFFSR_184 ( );
FILL FILL_1_DFFSR_184 ( );
FILL FILL_2_DFFSR_184 ( );
FILL FILL_3_DFFSR_184 ( );
FILL FILL_4_DFFSR_184 ( );
FILL FILL_5_DFFSR_184 ( );
FILL FILL_6_DFFSR_184 ( );
FILL FILL_7_DFFSR_184 ( );
FILL FILL_8_DFFSR_184 ( );
FILL FILL_9_DFFSR_184 ( );
FILL FILL_10_DFFSR_184 ( );
FILL FILL_11_DFFSR_184 ( );
FILL FILL_12_DFFSR_184 ( );
FILL FILL_13_DFFSR_184 ( );
FILL FILL_14_DFFSR_184 ( );
FILL FILL_15_DFFSR_184 ( );
FILL FILL_16_DFFSR_184 ( );
FILL FILL_17_DFFSR_184 ( );
FILL FILL_18_DFFSR_184 ( );
FILL FILL_19_DFFSR_184 ( );
FILL FILL_20_DFFSR_184 ( );
FILL FILL_21_DFFSR_184 ( );
FILL FILL_22_DFFSR_184 ( );
FILL FILL_23_DFFSR_184 ( );
FILL FILL_24_DFFSR_184 ( );
FILL FILL_25_DFFSR_184 ( );
FILL FILL_26_DFFSR_184 ( );
FILL FILL_27_DFFSR_184 ( );
FILL FILL_28_DFFSR_184 ( );
FILL FILL_29_DFFSR_184 ( );
FILL FILL_30_DFFSR_184 ( );
FILL FILL_31_DFFSR_184 ( );
FILL FILL_32_DFFSR_184 ( );
FILL FILL_33_DFFSR_184 ( );
FILL FILL_34_DFFSR_184 ( );
FILL FILL_35_DFFSR_184 ( );
FILL FILL_36_DFFSR_184 ( );
FILL FILL_37_DFFSR_184 ( );
FILL FILL_38_DFFSR_184 ( );
FILL FILL_39_DFFSR_184 ( );
FILL FILL_40_DFFSR_184 ( );
FILL FILL_41_DFFSR_184 ( );
FILL FILL_42_DFFSR_184 ( );
FILL FILL_43_DFFSR_184 ( );
FILL FILL_44_DFFSR_184 ( );
FILL FILL_45_DFFSR_184 ( );
FILL FILL_46_DFFSR_184 ( );
FILL FILL_47_DFFSR_184 ( );
FILL FILL_48_DFFSR_184 ( );
FILL FILL_49_DFFSR_184 ( );
FILL FILL_50_DFFSR_184 ( );
FILL FILL_0_CLKBUF1_6 ( );
FILL FILL_1_CLKBUF1_6 ( );
FILL FILL_2_CLKBUF1_6 ( );
FILL FILL_3_CLKBUF1_6 ( );
FILL FILL_4_CLKBUF1_6 ( );
FILL FILL_5_CLKBUF1_6 ( );
FILL FILL_6_CLKBUF1_6 ( );
FILL FILL_7_CLKBUF1_6 ( );
FILL FILL_8_CLKBUF1_6 ( );
FILL FILL_9_CLKBUF1_6 ( );
FILL FILL_10_CLKBUF1_6 ( );
FILL FILL_11_CLKBUF1_6 ( );
FILL FILL_12_CLKBUF1_6 ( );
FILL FILL_13_CLKBUF1_6 ( );
FILL FILL_14_CLKBUF1_6 ( );
FILL FILL_15_CLKBUF1_6 ( );
FILL FILL_16_CLKBUF1_6 ( );
FILL FILL_17_CLKBUF1_6 ( );
FILL FILL_18_CLKBUF1_6 ( );
FILL FILL_19_CLKBUF1_6 ( );
FILL FILL_20_CLKBUF1_6 ( );
FILL FILL_0_NAND3X1_183 ( );
FILL FILL_1_NAND3X1_183 ( );
FILL FILL_2_NAND3X1_183 ( );
FILL FILL_3_NAND3X1_183 ( );
FILL FILL_4_NAND3X1_183 ( );
FILL FILL_5_NAND3X1_183 ( );
FILL FILL_6_NAND3X1_183 ( );
FILL FILL_7_NAND3X1_183 ( );
FILL FILL_8_NAND3X1_183 ( );
FILL FILL_0_NAND3X1_180 ( );
FILL FILL_1_NAND3X1_180 ( );
FILL FILL_2_NAND3X1_180 ( );
FILL FILL_3_NAND3X1_180 ( );
FILL FILL_4_NAND3X1_180 ( );
FILL FILL_5_NAND3X1_180 ( );
FILL FILL_6_NAND3X1_180 ( );
FILL FILL_7_NAND3X1_180 ( );
FILL FILL_8_NAND3X1_180 ( );
FILL FILL_0_NAND2X1_73 ( );
FILL FILL_1_NAND2X1_73 ( );
FILL FILL_2_NAND2X1_73 ( );
FILL FILL_3_NAND2X1_73 ( );
FILL FILL_4_NAND2X1_73 ( );
FILL FILL_5_NAND2X1_73 ( );
FILL FILL_6_NAND2X1_73 ( );
FILL FILL_0_OAI22X1_49 ( );
FILL FILL_1_OAI22X1_49 ( );
FILL FILL_2_OAI22X1_49 ( );
FILL FILL_3_OAI22X1_49 ( );
FILL FILL_4_OAI22X1_49 ( );
FILL FILL_5_OAI22X1_49 ( );
FILL FILL_6_OAI22X1_49 ( );
FILL FILL_7_OAI22X1_49 ( );
FILL FILL_8_OAI22X1_49 ( );
FILL FILL_9_OAI22X1_49 ( );
FILL FILL_10_OAI22X1_49 ( );
FILL FILL_11_OAI22X1_49 ( );
FILL FILL_0_NAND3X1_156 ( );
FILL FILL_1_NAND3X1_156 ( );
FILL FILL_2_NAND3X1_156 ( );
FILL FILL_3_NAND3X1_156 ( );
FILL FILL_4_NAND3X1_156 ( );
FILL FILL_5_NAND3X1_156 ( );
FILL FILL_6_NAND3X1_156 ( );
FILL FILL_7_NAND3X1_156 ( );
FILL FILL_8_NAND3X1_156 ( );
FILL FILL_0_AOI22X1_18 ( );
FILL FILL_1_AOI22X1_18 ( );
FILL FILL_2_AOI22X1_18 ( );
FILL FILL_3_AOI22X1_18 ( );
FILL FILL_4_AOI22X1_18 ( );
FILL FILL_5_AOI22X1_18 ( );
FILL FILL_6_AOI22X1_18 ( );
FILL FILL_7_AOI22X1_18 ( );
FILL FILL_8_AOI22X1_18 ( );
FILL FILL_9_AOI22X1_18 ( );
FILL FILL_10_AOI22X1_18 ( );
FILL FILL_0_OAI21X1_38 ( );
FILL FILL_1_OAI21X1_38 ( );
FILL FILL_2_OAI21X1_38 ( );
FILL FILL_3_OAI21X1_38 ( );
FILL FILL_4_OAI21X1_38 ( );
FILL FILL_5_OAI21X1_38 ( );
FILL FILL_6_OAI21X1_38 ( );
FILL FILL_7_OAI21X1_38 ( );
FILL FILL_8_OAI21X1_38 ( );
FILL FILL_9_OAI21X1_38 ( );
FILL FILL_0_DFFPOSX1_40 ( );
FILL FILL_1_DFFPOSX1_40 ( );
FILL FILL_2_DFFPOSX1_40 ( );
FILL FILL_3_DFFPOSX1_40 ( );
FILL FILL_4_DFFPOSX1_40 ( );
FILL FILL_5_DFFPOSX1_40 ( );
FILL FILL_6_DFFPOSX1_40 ( );
FILL FILL_7_DFFPOSX1_40 ( );
FILL FILL_8_DFFPOSX1_40 ( );
FILL FILL_9_DFFPOSX1_40 ( );
FILL FILL_10_DFFPOSX1_40 ( );
FILL FILL_11_DFFPOSX1_40 ( );
FILL FILL_12_DFFPOSX1_40 ( );
FILL FILL_13_DFFPOSX1_40 ( );
FILL FILL_14_DFFPOSX1_40 ( );
FILL FILL_15_DFFPOSX1_40 ( );
FILL FILL_16_DFFPOSX1_40 ( );
FILL FILL_17_DFFPOSX1_40 ( );
FILL FILL_18_DFFPOSX1_40 ( );
FILL FILL_19_DFFPOSX1_40 ( );
FILL FILL_20_DFFPOSX1_40 ( );
FILL FILL_21_DFFPOSX1_40 ( );
FILL FILL_22_DFFPOSX1_40 ( );
FILL FILL_23_DFFPOSX1_40 ( );
FILL FILL_24_DFFPOSX1_40 ( );
FILL FILL_25_DFFPOSX1_40 ( );
FILL FILL_26_DFFPOSX1_40 ( );
FILL FILL_27_DFFPOSX1_40 ( );
FILL FILL_0_NAND2X1_167 ( );
FILL FILL_1_NAND2X1_167 ( );
FILL FILL_2_NAND2X1_167 ( );
FILL FILL_3_NAND2X1_167 ( );
FILL FILL_4_NAND2X1_167 ( );
FILL FILL_5_NAND2X1_167 ( );
FILL FILL_6_NAND2X1_167 ( );
FILL FILL_0_BUFX2_35 ( );
FILL FILL_1_BUFX2_35 ( );
FILL FILL_2_BUFX2_35 ( );
FILL FILL_3_BUFX2_35 ( );
FILL FILL_4_BUFX2_35 ( );
FILL FILL_5_BUFX2_35 ( );
FILL FILL_6_BUFX2_35 ( );
FILL FILL_0_INVX1_59 ( );
FILL FILL_1_INVX1_59 ( );
FILL FILL_2_INVX1_59 ( );
FILL FILL_3_INVX1_59 ( );
FILL FILL_4_INVX1_59 ( );
FILL FILL_0_OR2X2_1 ( );
FILL FILL_1_OR2X2_1 ( );
FILL FILL_2_OR2X2_1 ( );
FILL FILL_3_OR2X2_1 ( );
FILL FILL_4_OR2X2_1 ( );
FILL FILL_5_OR2X2_1 ( );
FILL FILL_6_OR2X2_1 ( );
FILL FILL_7_OR2X2_1 ( );
FILL FILL_8_OR2X2_1 ( );
FILL FILL_0_DFFPOSX1_45 ( );
FILL FILL_1_DFFPOSX1_45 ( );
FILL FILL_2_DFFPOSX1_45 ( );
FILL FILL_3_DFFPOSX1_45 ( );
FILL FILL_4_DFFPOSX1_45 ( );
FILL FILL_5_DFFPOSX1_45 ( );
FILL FILL_6_DFFPOSX1_45 ( );
FILL FILL_7_DFFPOSX1_45 ( );
FILL FILL_8_DFFPOSX1_45 ( );
FILL FILL_9_DFFPOSX1_45 ( );
FILL FILL_10_DFFPOSX1_45 ( );
FILL FILL_11_DFFPOSX1_45 ( );
FILL FILL_12_DFFPOSX1_45 ( );
FILL FILL_13_DFFPOSX1_45 ( );
FILL FILL_14_DFFPOSX1_45 ( );
FILL FILL_15_DFFPOSX1_45 ( );
FILL FILL_16_DFFPOSX1_45 ( );
FILL FILL_17_DFFPOSX1_45 ( );
FILL FILL_18_DFFPOSX1_45 ( );
FILL FILL_19_DFFPOSX1_45 ( );
FILL FILL_20_DFFPOSX1_45 ( );
FILL FILL_21_DFFPOSX1_45 ( );
FILL FILL_22_DFFPOSX1_45 ( );
FILL FILL_23_DFFPOSX1_45 ( );
FILL FILL_24_DFFPOSX1_45 ( );
FILL FILL_25_DFFPOSX1_45 ( );
FILL FILL_26_DFFPOSX1_45 ( );
FILL FILL_27_DFFPOSX1_45 ( );
FILL FILL_0_BUFX2_10 ( );
FILL FILL_1_BUFX2_10 ( );
FILL FILL_2_BUFX2_10 ( );
FILL FILL_3_BUFX2_10 ( );
FILL FILL_4_BUFX2_10 ( );
FILL FILL_5_BUFX2_10 ( );
FILL FILL_0_DFFSR_124 ( );
FILL FILL_1_DFFSR_124 ( );
FILL FILL_2_DFFSR_124 ( );
FILL FILL_3_DFFSR_124 ( );
FILL FILL_4_DFFSR_124 ( );
FILL FILL_5_DFFSR_124 ( );
FILL FILL_6_DFFSR_124 ( );
FILL FILL_7_DFFSR_124 ( );
FILL FILL_8_DFFSR_124 ( );
FILL FILL_9_DFFSR_124 ( );
FILL FILL_10_DFFSR_124 ( );
FILL FILL_11_DFFSR_124 ( );
FILL FILL_12_DFFSR_124 ( );
FILL FILL_13_DFFSR_124 ( );
FILL FILL_14_DFFSR_124 ( );
FILL FILL_15_DFFSR_124 ( );
FILL FILL_16_DFFSR_124 ( );
FILL FILL_17_DFFSR_124 ( );
FILL FILL_18_DFFSR_124 ( );
FILL FILL_19_DFFSR_124 ( );
FILL FILL_20_DFFSR_124 ( );
FILL FILL_21_DFFSR_124 ( );
FILL FILL_22_DFFSR_124 ( );
FILL FILL_23_DFFSR_124 ( );
FILL FILL_24_DFFSR_124 ( );
FILL FILL_25_DFFSR_124 ( );
FILL FILL_26_DFFSR_124 ( );
FILL FILL_27_DFFSR_124 ( );
FILL FILL_28_DFFSR_124 ( );
FILL FILL_29_DFFSR_124 ( );
FILL FILL_30_DFFSR_124 ( );
FILL FILL_31_DFFSR_124 ( );
FILL FILL_32_DFFSR_124 ( );
FILL FILL_33_DFFSR_124 ( );
FILL FILL_34_DFFSR_124 ( );
FILL FILL_35_DFFSR_124 ( );
FILL FILL_36_DFFSR_124 ( );
FILL FILL_37_DFFSR_124 ( );
FILL FILL_38_DFFSR_124 ( );
FILL FILL_39_DFFSR_124 ( );
FILL FILL_40_DFFSR_124 ( );
FILL FILL_41_DFFSR_124 ( );
FILL FILL_42_DFFSR_124 ( );
FILL FILL_43_DFFSR_124 ( );
FILL FILL_44_DFFSR_124 ( );
FILL FILL_45_DFFSR_124 ( );
FILL FILL_46_DFFSR_124 ( );
FILL FILL_47_DFFSR_124 ( );
FILL FILL_48_DFFSR_124 ( );
FILL FILL_49_DFFSR_124 ( );
FILL FILL_50_DFFSR_124 ( );
FILL FILL_0_INVX1_187 ( );
FILL FILL_1_INVX1_187 ( );
FILL FILL_2_INVX1_187 ( );
FILL FILL_3_INVX1_187 ( );
FILL FILL_4_INVX1_187 ( );
FILL FILL_0_INVX1_18 ( );
FILL FILL_1_INVX1_18 ( );
FILL FILL_2_INVX1_18 ( );
FILL FILL_3_INVX1_18 ( );
FILL FILL_0_XOR2X1_10 ( );
FILL FILL_1_XOR2X1_10 ( );
FILL FILL_2_XOR2X1_10 ( );
FILL FILL_3_XOR2X1_10 ( );
FILL FILL_4_XOR2X1_10 ( );
FILL FILL_5_XOR2X1_10 ( );
FILL FILL_6_XOR2X1_10 ( );
FILL FILL_7_XOR2X1_10 ( );
FILL FILL_8_XOR2X1_10 ( );
FILL FILL_9_XOR2X1_10 ( );
FILL FILL_10_XOR2X1_10 ( );
FILL FILL_11_XOR2X1_10 ( );
FILL FILL_12_XOR2X1_10 ( );
FILL FILL_13_XOR2X1_10 ( );
FILL FILL_14_XOR2X1_10 ( );
FILL FILL_15_XOR2X1_10 ( );
FILL FILL_0_NAND2X1_172 ( );
FILL FILL_1_NAND2X1_172 ( );
FILL FILL_2_NAND2X1_172 ( );
FILL FILL_3_NAND2X1_172 ( );
FILL FILL_4_NAND2X1_172 ( );
FILL FILL_5_NAND2X1_172 ( );
FILL FILL_6_NAND2X1_172 ( );
FILL FILL_0_DFFSR_89 ( );
FILL FILL_1_DFFSR_89 ( );
FILL FILL_2_DFFSR_89 ( );
FILL FILL_3_DFFSR_89 ( );
FILL FILL_4_DFFSR_89 ( );
FILL FILL_5_DFFSR_89 ( );
FILL FILL_6_DFFSR_89 ( );
FILL FILL_7_DFFSR_89 ( );
FILL FILL_8_DFFSR_89 ( );
FILL FILL_9_DFFSR_89 ( );
FILL FILL_10_DFFSR_89 ( );
FILL FILL_11_DFFSR_89 ( );
FILL FILL_12_DFFSR_89 ( );
FILL FILL_13_DFFSR_89 ( );
FILL FILL_14_DFFSR_89 ( );
FILL FILL_15_DFFSR_89 ( );
FILL FILL_16_DFFSR_89 ( );
FILL FILL_17_DFFSR_89 ( );
FILL FILL_18_DFFSR_89 ( );
FILL FILL_19_DFFSR_89 ( );
FILL FILL_20_DFFSR_89 ( );
FILL FILL_21_DFFSR_89 ( );
FILL FILL_22_DFFSR_89 ( );
FILL FILL_23_DFFSR_89 ( );
FILL FILL_24_DFFSR_89 ( );
FILL FILL_25_DFFSR_89 ( );
FILL FILL_26_DFFSR_89 ( );
FILL FILL_27_DFFSR_89 ( );
FILL FILL_28_DFFSR_89 ( );
FILL FILL_29_DFFSR_89 ( );
FILL FILL_30_DFFSR_89 ( );
FILL FILL_31_DFFSR_89 ( );
FILL FILL_32_DFFSR_89 ( );
FILL FILL_33_DFFSR_89 ( );
FILL FILL_34_DFFSR_89 ( );
FILL FILL_35_DFFSR_89 ( );
FILL FILL_36_DFFSR_89 ( );
FILL FILL_37_DFFSR_89 ( );
FILL FILL_38_DFFSR_89 ( );
FILL FILL_39_DFFSR_89 ( );
FILL FILL_40_DFFSR_89 ( );
FILL FILL_41_DFFSR_89 ( );
FILL FILL_42_DFFSR_89 ( );
FILL FILL_43_DFFSR_89 ( );
FILL FILL_44_DFFSR_89 ( );
FILL FILL_45_DFFSR_89 ( );
FILL FILL_46_DFFSR_89 ( );
FILL FILL_47_DFFSR_89 ( );
FILL FILL_48_DFFSR_89 ( );
FILL FILL_49_DFFSR_89 ( );
FILL FILL_50_DFFSR_89 ( );
FILL FILL_51_DFFSR_89 ( );
FILL FILL_0_AND2X2_22 ( );
FILL FILL_1_AND2X2_22 ( );
FILL FILL_2_AND2X2_22 ( );
FILL FILL_3_AND2X2_22 ( );
FILL FILL_4_AND2X2_22 ( );
FILL FILL_5_AND2X2_22 ( );
FILL FILL_6_AND2X2_22 ( );
FILL FILL_7_AND2X2_22 ( );
FILL FILL_8_AND2X2_22 ( );
FILL FILL_0_NAND3X1_90 ( );
FILL FILL_1_NAND3X1_90 ( );
FILL FILL_2_NAND3X1_90 ( );
FILL FILL_3_NAND3X1_90 ( );
FILL FILL_4_NAND3X1_90 ( );
FILL FILL_5_NAND3X1_90 ( );
FILL FILL_6_NAND3X1_90 ( );
FILL FILL_7_NAND3X1_90 ( );
FILL FILL_8_NAND3X1_90 ( );
FILL FILL_0_DFFSR_155 ( );
FILL FILL_1_DFFSR_155 ( );
FILL FILL_2_DFFSR_155 ( );
FILL FILL_3_DFFSR_155 ( );
FILL FILL_4_DFFSR_155 ( );
FILL FILL_5_DFFSR_155 ( );
FILL FILL_6_DFFSR_155 ( );
FILL FILL_7_DFFSR_155 ( );
FILL FILL_8_DFFSR_155 ( );
FILL FILL_9_DFFSR_155 ( );
FILL FILL_10_DFFSR_155 ( );
FILL FILL_11_DFFSR_155 ( );
FILL FILL_12_DFFSR_155 ( );
FILL FILL_13_DFFSR_155 ( );
FILL FILL_14_DFFSR_155 ( );
FILL FILL_15_DFFSR_155 ( );
FILL FILL_16_DFFSR_155 ( );
FILL FILL_17_DFFSR_155 ( );
FILL FILL_18_DFFSR_155 ( );
FILL FILL_19_DFFSR_155 ( );
FILL FILL_20_DFFSR_155 ( );
FILL FILL_21_DFFSR_155 ( );
FILL FILL_22_DFFSR_155 ( );
FILL FILL_23_DFFSR_155 ( );
FILL FILL_24_DFFSR_155 ( );
FILL FILL_25_DFFSR_155 ( );
FILL FILL_26_DFFSR_155 ( );
FILL FILL_27_DFFSR_155 ( );
FILL FILL_28_DFFSR_155 ( );
FILL FILL_29_DFFSR_155 ( );
FILL FILL_30_DFFSR_155 ( );
FILL FILL_31_DFFSR_155 ( );
FILL FILL_32_DFFSR_155 ( );
FILL FILL_33_DFFSR_155 ( );
FILL FILL_34_DFFSR_155 ( );
FILL FILL_35_DFFSR_155 ( );
FILL FILL_36_DFFSR_155 ( );
FILL FILL_37_DFFSR_155 ( );
FILL FILL_38_DFFSR_155 ( );
FILL FILL_39_DFFSR_155 ( );
FILL FILL_40_DFFSR_155 ( );
FILL FILL_41_DFFSR_155 ( );
FILL FILL_42_DFFSR_155 ( );
FILL FILL_43_DFFSR_155 ( );
FILL FILL_44_DFFSR_155 ( );
FILL FILL_45_DFFSR_155 ( );
FILL FILL_46_DFFSR_155 ( );
FILL FILL_47_DFFSR_155 ( );
FILL FILL_48_DFFSR_155 ( );
FILL FILL_49_DFFSR_155 ( );
FILL FILL_50_DFFSR_155 ( );
FILL FILL_51_DFFSR_155 ( );
FILL FILL_0_INVX1_102 ( );
FILL FILL_1_INVX1_102 ( );
FILL FILL_2_INVX1_102 ( );
FILL FILL_3_INVX1_102 ( );
FILL FILL_0_CLKBUF1_22 ( );
FILL FILL_1_CLKBUF1_22 ( );
FILL FILL_2_CLKBUF1_22 ( );
FILL FILL_3_CLKBUF1_22 ( );
FILL FILL_4_CLKBUF1_22 ( );
FILL FILL_5_CLKBUF1_22 ( );
FILL FILL_6_CLKBUF1_22 ( );
FILL FILL_7_CLKBUF1_22 ( );
FILL FILL_8_CLKBUF1_22 ( );
FILL FILL_9_CLKBUF1_22 ( );
FILL FILL_10_CLKBUF1_22 ( );
FILL FILL_11_CLKBUF1_22 ( );
FILL FILL_12_CLKBUF1_22 ( );
FILL FILL_13_CLKBUF1_22 ( );
FILL FILL_14_CLKBUF1_22 ( );
FILL FILL_15_CLKBUF1_22 ( );
FILL FILL_16_CLKBUF1_22 ( );
FILL FILL_17_CLKBUF1_22 ( );
FILL FILL_18_CLKBUF1_22 ( );
FILL FILL_19_CLKBUF1_22 ( );
FILL FILL_20_CLKBUF1_22 ( );
FILL FILL_0_NAND3X1_98 ( );
FILL FILL_1_NAND3X1_98 ( );
FILL FILL_2_NAND3X1_98 ( );
FILL FILL_3_NAND3X1_98 ( );
FILL FILL_4_NAND3X1_98 ( );
FILL FILL_5_NAND3X1_98 ( );
FILL FILL_6_NAND3X1_98 ( );
FILL FILL_7_NAND3X1_98 ( );
FILL FILL_8_NAND3X1_98 ( );
FILL FILL_0_AND2X2_23 ( );
FILL FILL_1_AND2X2_23 ( );
FILL FILL_2_AND2X2_23 ( );
FILL FILL_3_AND2X2_23 ( );
FILL FILL_4_AND2X2_23 ( );
FILL FILL_5_AND2X2_23 ( );
FILL FILL_6_AND2X2_23 ( );
FILL FILL_7_AND2X2_23 ( );
FILL FILL_8_AND2X2_23 ( );
FILL FILL_9_AND2X2_23 ( );
FILL FILL_0_OAI22X1_46 ( );
FILL FILL_1_OAI22X1_46 ( );
FILL FILL_2_OAI22X1_46 ( );
FILL FILL_3_OAI22X1_46 ( );
FILL FILL_4_OAI22X1_46 ( );
FILL FILL_5_OAI22X1_46 ( );
FILL FILL_6_OAI22X1_46 ( );
FILL FILL_7_OAI22X1_46 ( );
FILL FILL_8_OAI22X1_46 ( );
FILL FILL_9_OAI22X1_46 ( );
FILL FILL_10_OAI22X1_46 ( );
FILL FILL_0_INVX1_111 ( );
FILL FILL_1_INVX1_111 ( );
FILL FILL_2_INVX1_111 ( );
FILL FILL_3_INVX1_111 ( );
FILL FILL_4_INVX1_111 ( );
FILL FILL_0_DFFSR_229 ( );
FILL FILL_1_DFFSR_229 ( );
FILL FILL_2_DFFSR_229 ( );
FILL FILL_3_DFFSR_229 ( );
FILL FILL_4_DFFSR_229 ( );
FILL FILL_5_DFFSR_229 ( );
FILL FILL_6_DFFSR_229 ( );
FILL FILL_7_DFFSR_229 ( );
FILL FILL_8_DFFSR_229 ( );
FILL FILL_9_DFFSR_229 ( );
FILL FILL_10_DFFSR_229 ( );
FILL FILL_11_DFFSR_229 ( );
FILL FILL_12_DFFSR_229 ( );
FILL FILL_13_DFFSR_229 ( );
FILL FILL_14_DFFSR_229 ( );
FILL FILL_15_DFFSR_229 ( );
FILL FILL_16_DFFSR_229 ( );
FILL FILL_17_DFFSR_229 ( );
FILL FILL_18_DFFSR_229 ( );
FILL FILL_19_DFFSR_229 ( );
FILL FILL_20_DFFSR_229 ( );
FILL FILL_21_DFFSR_229 ( );
FILL FILL_22_DFFSR_229 ( );
FILL FILL_23_DFFSR_229 ( );
FILL FILL_24_DFFSR_229 ( );
FILL FILL_25_DFFSR_229 ( );
FILL FILL_26_DFFSR_229 ( );
FILL FILL_27_DFFSR_229 ( );
FILL FILL_28_DFFSR_229 ( );
FILL FILL_29_DFFSR_229 ( );
FILL FILL_30_DFFSR_229 ( );
FILL FILL_31_DFFSR_229 ( );
FILL FILL_32_DFFSR_229 ( );
FILL FILL_33_DFFSR_229 ( );
FILL FILL_34_DFFSR_229 ( );
FILL FILL_35_DFFSR_229 ( );
FILL FILL_36_DFFSR_229 ( );
FILL FILL_37_DFFSR_229 ( );
FILL FILL_38_DFFSR_229 ( );
FILL FILL_39_DFFSR_229 ( );
FILL FILL_40_DFFSR_229 ( );
FILL FILL_41_DFFSR_229 ( );
FILL FILL_42_DFFSR_229 ( );
FILL FILL_43_DFFSR_229 ( );
FILL FILL_44_DFFSR_229 ( );
FILL FILL_45_DFFSR_229 ( );
FILL FILL_46_DFFSR_229 ( );
FILL FILL_47_DFFSR_229 ( );
FILL FILL_48_DFFSR_229 ( );
FILL FILL_49_DFFSR_229 ( );
FILL FILL_50_DFFSR_229 ( );
FILL FILL_51_DFFSR_229 ( );
FILL FILL_0_AND2X2_38 ( );
FILL FILL_1_AND2X2_38 ( );
FILL FILL_2_AND2X2_38 ( );
FILL FILL_3_AND2X2_38 ( );
FILL FILL_4_AND2X2_38 ( );
FILL FILL_5_AND2X2_38 ( );
FILL FILL_6_AND2X2_38 ( );
FILL FILL_7_AND2X2_38 ( );
FILL FILL_8_AND2X2_38 ( );
FILL FILL_9_AND2X2_38 ( );
FILL FILL_0_NAND2X1_72 ( );
FILL FILL_1_NAND2X1_72 ( );
FILL FILL_2_NAND2X1_72 ( );
FILL FILL_3_NAND2X1_72 ( );
FILL FILL_4_NAND2X1_72 ( );
FILL FILL_5_NAND2X1_72 ( );
FILL FILL_6_NAND2X1_72 ( );
FILL FILL_0_NAND3X1_177 ( );
FILL FILL_1_NAND3X1_177 ( );
FILL FILL_2_NAND3X1_177 ( );
FILL FILL_3_NAND3X1_177 ( );
FILL FILL_4_NAND3X1_177 ( );
FILL FILL_5_NAND3X1_177 ( );
FILL FILL_6_NAND3X1_177 ( );
FILL FILL_7_NAND3X1_177 ( );
FILL FILL_8_NAND3X1_177 ( );
FILL FILL_0_AOI22X1_21 ( );
FILL FILL_1_AOI22X1_21 ( );
FILL FILL_2_AOI22X1_21 ( );
FILL FILL_3_AOI22X1_21 ( );
FILL FILL_4_AOI22X1_21 ( );
FILL FILL_5_AOI22X1_21 ( );
FILL FILL_6_AOI22X1_21 ( );
FILL FILL_7_AOI22X1_21 ( );
FILL FILL_8_AOI22X1_21 ( );
FILL FILL_9_AOI22X1_21 ( );
FILL FILL_10_AOI22X1_21 ( );
FILL FILL_0_NAND2X1_74 ( );
FILL FILL_1_NAND2X1_74 ( );
FILL FILL_2_NAND2X1_74 ( );
FILL FILL_3_NAND2X1_74 ( );
FILL FILL_4_NAND2X1_74 ( );
FILL FILL_5_NAND2X1_74 ( );
FILL FILL_6_NAND2X1_74 ( );
FILL FILL_0_NAND3X1_158 ( );
FILL FILL_1_NAND3X1_158 ( );
FILL FILL_2_NAND3X1_158 ( );
FILL FILL_3_NAND3X1_158 ( );
FILL FILL_4_NAND3X1_158 ( );
FILL FILL_5_NAND3X1_158 ( );
FILL FILL_6_NAND3X1_158 ( );
FILL FILL_7_NAND3X1_158 ( );
FILL FILL_8_NAND3X1_158 ( );
FILL FILL_0_OAI21X1_32 ( );
FILL FILL_1_OAI21X1_32 ( );
FILL FILL_2_OAI21X1_32 ( );
FILL FILL_3_OAI21X1_32 ( );
FILL FILL_4_OAI21X1_32 ( );
FILL FILL_5_OAI21X1_32 ( );
FILL FILL_6_OAI21X1_32 ( );
FILL FILL_7_OAI21X1_32 ( );
FILL FILL_8_OAI21X1_32 ( );
FILL FILL_9_OAI21X1_32 ( );
FILL FILL_0_NAND3X1_144 ( );
FILL FILL_1_NAND3X1_144 ( );
FILL FILL_2_NAND3X1_144 ( );
FILL FILL_3_NAND3X1_144 ( );
FILL FILL_4_NAND3X1_144 ( );
FILL FILL_5_NAND3X1_144 ( );
FILL FILL_6_NAND3X1_144 ( );
FILL FILL_7_NAND3X1_144 ( );
FILL FILL_8_NAND3X1_144 ( );
FILL FILL_0_NAND2X1_67 ( );
FILL FILL_1_NAND2X1_67 ( );
FILL FILL_2_NAND2X1_67 ( );
FILL FILL_3_NAND2X1_67 ( );
FILL FILL_4_NAND2X1_67 ( );
FILL FILL_5_NAND2X1_67 ( );
FILL FILL_6_NAND2X1_67 ( );
FILL FILL_0_AND2X2_34 ( );
FILL FILL_1_AND2X2_34 ( );
FILL FILL_2_AND2X2_34 ( );
FILL FILL_3_AND2X2_34 ( );
FILL FILL_4_AND2X2_34 ( );
FILL FILL_5_AND2X2_34 ( );
FILL FILL_6_AND2X2_34 ( );
FILL FILL_7_AND2X2_34 ( );
FILL FILL_8_AND2X2_34 ( );
FILL FILL_9_AND2X2_34 ( );
FILL FILL_0_OAI21X1_96 ( );
FILL FILL_1_OAI21X1_96 ( );
FILL FILL_2_OAI21X1_96 ( );
FILL FILL_3_OAI21X1_96 ( );
FILL FILL_4_OAI21X1_96 ( );
FILL FILL_5_OAI21X1_96 ( );
FILL FILL_6_OAI21X1_96 ( );
FILL FILL_7_OAI21X1_96 ( );
FILL FILL_8_OAI21X1_96 ( );
FILL FILL_9_OAI21X1_96 ( );
FILL FILL_0_NAND2X1_63 ( );
FILL FILL_1_NAND2X1_63 ( );
FILL FILL_2_NAND2X1_63 ( );
FILL FILL_3_NAND2X1_63 ( );
FILL FILL_4_NAND2X1_63 ( );
FILL FILL_5_NAND2X1_63 ( );
FILL FILL_6_NAND2X1_63 ( );
FILL FILL_0_AOI21X1_54 ( );
FILL FILL_1_AOI21X1_54 ( );
FILL FILL_2_AOI21X1_54 ( );
FILL FILL_3_AOI21X1_54 ( );
FILL FILL_4_AOI21X1_54 ( );
FILL FILL_5_AOI21X1_54 ( );
FILL FILL_6_AOI21X1_54 ( );
FILL FILL_7_AOI21X1_54 ( );
FILL FILL_8_AOI21X1_54 ( );
FILL FILL_0_NAND2X1_156 ( );
FILL FILL_1_NAND2X1_156 ( );
FILL FILL_2_NAND2X1_156 ( );
FILL FILL_3_NAND2X1_156 ( );
FILL FILL_4_NAND2X1_156 ( );
FILL FILL_5_NAND2X1_156 ( );
FILL FILL_6_NAND2X1_156 ( );
FILL FILL_0_AOI21X1_61 ( );
FILL FILL_1_AOI21X1_61 ( );
FILL FILL_2_AOI21X1_61 ( );
FILL FILL_3_AOI21X1_61 ( );
FILL FILL_4_AOI21X1_61 ( );
FILL FILL_5_AOI21X1_61 ( );
FILL FILL_6_AOI21X1_61 ( );
FILL FILL_7_AOI21X1_61 ( );
FILL FILL_8_AOI21X1_61 ( );
FILL FILL_0_NOR2X1_64 ( );
FILL FILL_1_NOR2X1_64 ( );
FILL FILL_2_NOR2X1_64 ( );
FILL FILL_3_NOR2X1_64 ( );
FILL FILL_4_NOR2X1_64 ( );
FILL FILL_5_NOR2X1_64 ( );
FILL FILL_6_NOR2X1_64 ( );
FILL FILL_0_OAI21X1_21 ( );
FILL FILL_1_OAI21X1_21 ( );
FILL FILL_2_OAI21X1_21 ( );
FILL FILL_3_OAI21X1_21 ( );
FILL FILL_4_OAI21X1_21 ( );
FILL FILL_5_OAI21X1_21 ( );
FILL FILL_6_OAI21X1_21 ( );
FILL FILL_7_OAI21X1_21 ( );
FILL FILL_8_OAI21X1_21 ( );
FILL FILL_9_OAI21X1_21 ( );
FILL FILL_0_NAND2X1_56 ( );
FILL FILL_1_NAND2X1_56 ( );
FILL FILL_2_NAND2X1_56 ( );
FILL FILL_3_NAND2X1_56 ( );
FILL FILL_4_NAND2X1_56 ( );
FILL FILL_5_NAND2X1_56 ( );
FILL FILL_6_NAND2X1_56 ( );
FILL FILL_0_BUFX2_9 ( );
FILL FILL_1_BUFX2_9 ( );
FILL FILL_2_BUFX2_9 ( );
FILL FILL_3_BUFX2_9 ( );
FILL FILL_4_BUFX2_9 ( );
FILL FILL_5_BUFX2_9 ( );
FILL FILL_6_BUFX2_9 ( );
FILL FILL_7_BUFX2_9 ( );
FILL FILL_0_AOI21X1_64 ( );
FILL FILL_1_AOI21X1_64 ( );
FILL FILL_2_AOI21X1_64 ( );
FILL FILL_3_AOI21X1_64 ( );
FILL FILL_4_AOI21X1_64 ( );
FILL FILL_5_AOI21X1_64 ( );
FILL FILL_6_AOI21X1_64 ( );
FILL FILL_7_AOI21X1_64 ( );
FILL FILL_8_AOI21X1_64 ( );
FILL FILL_0_OAI21X1_114 ( );
FILL FILL_1_OAI21X1_114 ( );
FILL FILL_2_OAI21X1_114 ( );
FILL FILL_3_OAI21X1_114 ( );
FILL FILL_4_OAI21X1_114 ( );
FILL FILL_5_OAI21X1_114 ( );
FILL FILL_6_OAI21X1_114 ( );
FILL FILL_7_OAI21X1_114 ( );
FILL FILL_8_OAI21X1_114 ( );
FILL FILL_9_OAI21X1_114 ( );
FILL FILL_0_NAND2X1_54 ( );
FILL FILL_1_NAND2X1_54 ( );
FILL FILL_2_NAND2X1_54 ( );
FILL FILL_3_NAND2X1_54 ( );
FILL FILL_4_NAND2X1_54 ( );
FILL FILL_5_NAND2X1_54 ( );
FILL FILL_6_NAND2X1_54 ( );
FILL FILL_0_OAI22X1_16 ( );
FILL FILL_1_OAI22X1_16 ( );
FILL FILL_2_OAI22X1_16 ( );
FILL FILL_3_OAI22X1_16 ( );
FILL FILL_4_OAI22X1_16 ( );
FILL FILL_5_OAI22X1_16 ( );
FILL FILL_6_OAI22X1_16 ( );
FILL FILL_7_OAI22X1_16 ( );
FILL FILL_8_OAI22X1_16 ( );
FILL FILL_9_OAI22X1_16 ( );
FILL FILL_10_OAI22X1_16 ( );
FILL FILL_11_OAI22X1_16 ( );
FILL FILL_0_INVX1_17 ( );
FILL FILL_1_INVX1_17 ( );
FILL FILL_2_INVX1_17 ( );
FILL FILL_3_INVX1_17 ( );
FILL FILL_4_INVX1_17 ( );
FILL FILL_0_OAI22X1_7 ( );
FILL FILL_1_OAI22X1_7 ( );
FILL FILL_2_OAI22X1_7 ( );
FILL FILL_3_OAI22X1_7 ( );
FILL FILL_4_OAI22X1_7 ( );
FILL FILL_5_OAI22X1_7 ( );
FILL FILL_6_OAI22X1_7 ( );
FILL FILL_7_OAI22X1_7 ( );
FILL FILL_8_OAI22X1_7 ( );
FILL FILL_9_OAI22X1_7 ( );
FILL FILL_10_OAI22X1_7 ( );
FILL FILL_11_OAI22X1_7 ( );
FILL FILL_0_OAI21X1_111 ( );
FILL FILL_1_OAI21X1_111 ( );
FILL FILL_2_OAI21X1_111 ( );
FILL FILL_3_OAI21X1_111 ( );
FILL FILL_4_OAI21X1_111 ( );
FILL FILL_5_OAI21X1_111 ( );
FILL FILL_6_OAI21X1_111 ( );
FILL FILL_7_OAI21X1_111 ( );
FILL FILL_8_OAI21X1_111 ( );
FILL FILL_9_OAI21X1_111 ( );
FILL FILL_0_DFFSR_59 ( );
FILL FILL_1_DFFSR_59 ( );
FILL FILL_2_DFFSR_59 ( );
FILL FILL_3_DFFSR_59 ( );
FILL FILL_4_DFFSR_59 ( );
FILL FILL_5_DFFSR_59 ( );
FILL FILL_6_DFFSR_59 ( );
FILL FILL_7_DFFSR_59 ( );
FILL FILL_8_DFFSR_59 ( );
FILL FILL_9_DFFSR_59 ( );
FILL FILL_10_DFFSR_59 ( );
FILL FILL_11_DFFSR_59 ( );
FILL FILL_12_DFFSR_59 ( );
FILL FILL_13_DFFSR_59 ( );
FILL FILL_14_DFFSR_59 ( );
FILL FILL_15_DFFSR_59 ( );
FILL FILL_16_DFFSR_59 ( );
FILL FILL_17_DFFSR_59 ( );
FILL FILL_18_DFFSR_59 ( );
FILL FILL_19_DFFSR_59 ( );
FILL FILL_20_DFFSR_59 ( );
FILL FILL_21_DFFSR_59 ( );
FILL FILL_22_DFFSR_59 ( );
FILL FILL_23_DFFSR_59 ( );
FILL FILL_24_DFFSR_59 ( );
FILL FILL_25_DFFSR_59 ( );
FILL FILL_26_DFFSR_59 ( );
FILL FILL_27_DFFSR_59 ( );
FILL FILL_28_DFFSR_59 ( );
FILL FILL_29_DFFSR_59 ( );
FILL FILL_30_DFFSR_59 ( );
FILL FILL_31_DFFSR_59 ( );
FILL FILL_32_DFFSR_59 ( );
FILL FILL_33_DFFSR_59 ( );
FILL FILL_34_DFFSR_59 ( );
FILL FILL_35_DFFSR_59 ( );
FILL FILL_36_DFFSR_59 ( );
FILL FILL_37_DFFSR_59 ( );
FILL FILL_38_DFFSR_59 ( );
FILL FILL_39_DFFSR_59 ( );
FILL FILL_40_DFFSR_59 ( );
FILL FILL_41_DFFSR_59 ( );
FILL FILL_42_DFFSR_59 ( );
FILL FILL_43_DFFSR_59 ( );
FILL FILL_44_DFFSR_59 ( );
FILL FILL_45_DFFSR_59 ( );
FILL FILL_46_DFFSR_59 ( );
FILL FILL_47_DFFSR_59 ( );
FILL FILL_48_DFFSR_59 ( );
FILL FILL_49_DFFSR_59 ( );
FILL FILL_50_DFFSR_59 ( );
FILL FILL_0_BUFX2_48 ( );
FILL FILL_1_BUFX2_48 ( );
FILL FILL_2_BUFX2_48 ( );
FILL FILL_3_BUFX2_48 ( );
FILL FILL_4_BUFX2_48 ( );
FILL FILL_5_BUFX2_48 ( );
FILL FILL_6_BUFX2_48 ( );
FILL FILL_0_NAND3X1_131 ( );
FILL FILL_1_NAND3X1_131 ( );
FILL FILL_2_NAND3X1_131 ( );
FILL FILL_3_NAND3X1_131 ( );
FILL FILL_4_NAND3X1_131 ( );
FILL FILL_5_NAND3X1_131 ( );
FILL FILL_6_NAND3X1_131 ( );
FILL FILL_7_NAND3X1_131 ( );
FILL FILL_8_NAND3X1_131 ( );
FILL FILL_0_INVX1_125 ( );
FILL FILL_1_INVX1_125 ( );
FILL FILL_2_INVX1_125 ( );
FILL FILL_3_INVX1_125 ( );
FILL FILL_4_INVX1_125 ( );
FILL FILL_0_NAND3X1_91 ( );
FILL FILL_1_NAND3X1_91 ( );
FILL FILL_2_NAND3X1_91 ( );
FILL FILL_3_NAND3X1_91 ( );
FILL FILL_4_NAND3X1_91 ( );
FILL FILL_5_NAND3X1_91 ( );
FILL FILL_6_NAND3X1_91 ( );
FILL FILL_7_NAND3X1_91 ( );
FILL FILL_8_NAND3X1_91 ( );
FILL FILL_9_NAND3X1_91 ( );
FILL FILL_0_BUFX2_93 ( );
FILL FILL_1_BUFX2_93 ( );
FILL FILL_2_BUFX2_93 ( );
FILL FILL_3_BUFX2_93 ( );
FILL FILL_4_BUFX2_93 ( );
FILL FILL_5_BUFX2_93 ( );
FILL FILL_6_BUFX2_93 ( );
FILL FILL_0_NAND2X1_28 ( );
FILL FILL_1_NAND2X1_28 ( );
FILL FILL_2_NAND2X1_28 ( );
FILL FILL_3_NAND2X1_28 ( );
FILL FILL_4_NAND2X1_28 ( );
FILL FILL_5_NAND2X1_28 ( );
FILL FILL_6_NAND2X1_28 ( );
FILL FILL_0_DFFSR_166 ( );
FILL FILL_1_DFFSR_166 ( );
FILL FILL_2_DFFSR_166 ( );
FILL FILL_3_DFFSR_166 ( );
FILL FILL_4_DFFSR_166 ( );
FILL FILL_5_DFFSR_166 ( );
FILL FILL_6_DFFSR_166 ( );
FILL FILL_7_DFFSR_166 ( );
FILL FILL_8_DFFSR_166 ( );
FILL FILL_9_DFFSR_166 ( );
FILL FILL_10_DFFSR_166 ( );
FILL FILL_11_DFFSR_166 ( );
FILL FILL_12_DFFSR_166 ( );
FILL FILL_13_DFFSR_166 ( );
FILL FILL_14_DFFSR_166 ( );
FILL FILL_15_DFFSR_166 ( );
FILL FILL_16_DFFSR_166 ( );
FILL FILL_17_DFFSR_166 ( );
FILL FILL_18_DFFSR_166 ( );
FILL FILL_19_DFFSR_166 ( );
FILL FILL_20_DFFSR_166 ( );
FILL FILL_21_DFFSR_166 ( );
FILL FILL_22_DFFSR_166 ( );
FILL FILL_23_DFFSR_166 ( );
FILL FILL_24_DFFSR_166 ( );
FILL FILL_25_DFFSR_166 ( );
FILL FILL_26_DFFSR_166 ( );
FILL FILL_27_DFFSR_166 ( );
FILL FILL_28_DFFSR_166 ( );
FILL FILL_29_DFFSR_166 ( );
FILL FILL_30_DFFSR_166 ( );
FILL FILL_31_DFFSR_166 ( );
FILL FILL_32_DFFSR_166 ( );
FILL FILL_33_DFFSR_166 ( );
FILL FILL_34_DFFSR_166 ( );
FILL FILL_35_DFFSR_166 ( );
FILL FILL_36_DFFSR_166 ( );
FILL FILL_37_DFFSR_166 ( );
FILL FILL_38_DFFSR_166 ( );
FILL FILL_39_DFFSR_166 ( );
FILL FILL_40_DFFSR_166 ( );
FILL FILL_41_DFFSR_166 ( );
FILL FILL_42_DFFSR_166 ( );
FILL FILL_43_DFFSR_166 ( );
FILL FILL_44_DFFSR_166 ( );
FILL FILL_45_DFFSR_166 ( );
FILL FILL_46_DFFSR_166 ( );
FILL FILL_47_DFFSR_166 ( );
FILL FILL_48_DFFSR_166 ( );
FILL FILL_49_DFFSR_166 ( );
FILL FILL_50_DFFSR_166 ( );
FILL FILL_0_AND2X2_18 ( );
FILL FILL_1_AND2X2_18 ( );
FILL FILL_2_AND2X2_18 ( );
FILL FILL_3_AND2X2_18 ( );
FILL FILL_4_AND2X2_18 ( );
FILL FILL_5_AND2X2_18 ( );
FILL FILL_6_AND2X2_18 ( );
FILL FILL_7_AND2X2_18 ( );
FILL FILL_8_AND2X2_18 ( );
FILL FILL_0_BUFX2_5 ( );
FILL FILL_1_BUFX2_5 ( );
FILL FILL_2_BUFX2_5 ( );
FILL FILL_3_BUFX2_5 ( );
FILL FILL_4_BUFX2_5 ( );
FILL FILL_5_BUFX2_5 ( );
FILL FILL_6_BUFX2_5 ( );
FILL FILL_0_BUFX2_61 ( );
FILL FILL_1_BUFX2_61 ( );
FILL FILL_2_BUFX2_61 ( );
FILL FILL_3_BUFX2_61 ( );
FILL FILL_4_BUFX2_61 ( );
FILL FILL_5_BUFX2_61 ( );
FILL FILL_6_BUFX2_61 ( );
FILL FILL_0_NOR2X1_49 ( );
FILL FILL_1_NOR2X1_49 ( );
FILL FILL_2_NOR2X1_49 ( );
FILL FILL_3_NOR2X1_49 ( );
FILL FILL_4_NOR2X1_49 ( );
FILL FILL_5_NOR2X1_49 ( );
FILL FILL_6_NOR2X1_49 ( );
FILL FILL_0_NAND3X1_100 ( );
FILL FILL_1_NAND3X1_100 ( );
FILL FILL_2_NAND3X1_100 ( );
FILL FILL_3_NAND3X1_100 ( );
FILL FILL_4_NAND3X1_100 ( );
FILL FILL_5_NAND3X1_100 ( );
FILL FILL_6_NAND3X1_100 ( );
FILL FILL_7_NAND3X1_100 ( );
FILL FILL_8_NAND3X1_100 ( );
FILL FILL_0_NOR2X1_56 ( );
FILL FILL_1_NOR2X1_56 ( );
FILL FILL_2_NOR2X1_56 ( );
FILL FILL_3_NOR2X1_56 ( );
FILL FILL_4_NOR2X1_56 ( );
FILL FILL_5_NOR2X1_56 ( );
FILL FILL_6_NOR2X1_56 ( );
FILL FILL_0_NAND3X1_97 ( );
FILL FILL_1_NAND3X1_97 ( );
FILL FILL_2_NAND3X1_97 ( );
FILL FILL_3_NAND3X1_97 ( );
FILL FILL_4_NAND3X1_97 ( );
FILL FILL_5_NAND3X1_97 ( );
FILL FILL_6_NAND3X1_97 ( );
FILL FILL_7_NAND3X1_97 ( );
FILL FILL_8_NAND3X1_97 ( );
FILL FILL_9_NAND3X1_97 ( );
FILL FILL_0_DFFSR_221 ( );
FILL FILL_1_DFFSR_221 ( );
FILL FILL_2_DFFSR_221 ( );
FILL FILL_3_DFFSR_221 ( );
FILL FILL_4_DFFSR_221 ( );
FILL FILL_5_DFFSR_221 ( );
FILL FILL_6_DFFSR_221 ( );
FILL FILL_7_DFFSR_221 ( );
FILL FILL_8_DFFSR_221 ( );
FILL FILL_9_DFFSR_221 ( );
FILL FILL_10_DFFSR_221 ( );
FILL FILL_11_DFFSR_221 ( );
FILL FILL_12_DFFSR_221 ( );
FILL FILL_13_DFFSR_221 ( );
FILL FILL_14_DFFSR_221 ( );
FILL FILL_15_DFFSR_221 ( );
FILL FILL_16_DFFSR_221 ( );
FILL FILL_17_DFFSR_221 ( );
FILL FILL_18_DFFSR_221 ( );
FILL FILL_19_DFFSR_221 ( );
FILL FILL_20_DFFSR_221 ( );
FILL FILL_21_DFFSR_221 ( );
FILL FILL_22_DFFSR_221 ( );
FILL FILL_23_DFFSR_221 ( );
FILL FILL_24_DFFSR_221 ( );
FILL FILL_25_DFFSR_221 ( );
FILL FILL_26_DFFSR_221 ( );
FILL FILL_27_DFFSR_221 ( );
FILL FILL_28_DFFSR_221 ( );
FILL FILL_29_DFFSR_221 ( );
FILL FILL_30_DFFSR_221 ( );
FILL FILL_31_DFFSR_221 ( );
FILL FILL_32_DFFSR_221 ( );
FILL FILL_33_DFFSR_221 ( );
FILL FILL_34_DFFSR_221 ( );
FILL FILL_35_DFFSR_221 ( );
FILL FILL_36_DFFSR_221 ( );
FILL FILL_37_DFFSR_221 ( );
FILL FILL_38_DFFSR_221 ( );
FILL FILL_39_DFFSR_221 ( );
FILL FILL_40_DFFSR_221 ( );
FILL FILL_41_DFFSR_221 ( );
FILL FILL_42_DFFSR_221 ( );
FILL FILL_43_DFFSR_221 ( );
FILL FILL_44_DFFSR_221 ( );
FILL FILL_45_DFFSR_221 ( );
FILL FILL_46_DFFSR_221 ( );
FILL FILL_47_DFFSR_221 ( );
FILL FILL_48_DFFSR_221 ( );
FILL FILL_49_DFFSR_221 ( );
FILL FILL_50_DFFSR_221 ( );
FILL FILL_0_AOI21X1_28 ( );
FILL FILL_1_AOI21X1_28 ( );
FILL FILL_2_AOI21X1_28 ( );
FILL FILL_3_AOI21X1_28 ( );
FILL FILL_4_AOI21X1_28 ( );
FILL FILL_5_AOI21X1_28 ( );
FILL FILL_6_AOI21X1_28 ( );
FILL FILL_7_AOI21X1_28 ( );
FILL FILL_8_AOI21X1_28 ( );
FILL FILL_0_NAND2X1_103 ( );
FILL FILL_1_NAND2X1_103 ( );
FILL FILL_2_NAND2X1_103 ( );
FILL FILL_3_NAND2X1_103 ( );
FILL FILL_4_NAND2X1_103 ( );
FILL FILL_5_NAND2X1_103 ( );
FILL FILL_6_NAND2X1_103 ( );
FILL FILL_0_AND2X2_32 ( );
FILL FILL_1_AND2X2_32 ( );
FILL FILL_2_AND2X2_32 ( );
FILL FILL_3_AND2X2_32 ( );
FILL FILL_4_AND2X2_32 ( );
FILL FILL_5_AND2X2_32 ( );
FILL FILL_6_AND2X2_32 ( );
FILL FILL_7_AND2X2_32 ( );
FILL FILL_8_AND2X2_32 ( );
FILL FILL_0_OAI21X1_31 ( );
FILL FILL_1_OAI21X1_31 ( );
FILL FILL_2_OAI21X1_31 ( );
FILL FILL_3_OAI21X1_31 ( );
FILL FILL_4_OAI21X1_31 ( );
FILL FILL_5_OAI21X1_31 ( );
FILL FILL_6_OAI21X1_31 ( );
FILL FILL_7_OAI21X1_31 ( );
FILL FILL_8_OAI21X1_31 ( );
FILL FILL_0_NAND3X1_161 ( );
FILL FILL_1_NAND3X1_161 ( );
FILL FILL_2_NAND3X1_161 ( );
FILL FILL_3_NAND3X1_161 ( );
FILL FILL_4_NAND3X1_161 ( );
FILL FILL_5_NAND3X1_161 ( );
FILL FILL_6_NAND3X1_161 ( );
FILL FILL_7_NAND3X1_161 ( );
FILL FILL_8_NAND3X1_161 ( );
FILL FILL_9_NAND3X1_161 ( );
FILL FILL_0_NAND2X1_77 ( );
FILL FILL_1_NAND2X1_77 ( );
FILL FILL_2_NAND2X1_77 ( );
FILL FILL_3_NAND2X1_77 ( );
FILL FILL_4_NAND2X1_77 ( );
FILL FILL_5_NAND2X1_77 ( );
FILL FILL_6_NAND2X1_77 ( );
FILL FILL_0_NAND2X1_78 ( );
FILL FILL_1_NAND2X1_78 ( );
FILL FILL_2_NAND2X1_78 ( );
FILL FILL_3_NAND2X1_78 ( );
FILL FILL_4_NAND2X1_78 ( );
FILL FILL_5_NAND2X1_78 ( );
FILL FILL_6_NAND2X1_78 ( );
FILL FILL_0_NAND2X1_68 ( );
FILL FILL_1_NAND2X1_68 ( );
FILL FILL_2_NAND2X1_68 ( );
FILL FILL_3_NAND2X1_68 ( );
FILL FILL_4_NAND2X1_68 ( );
FILL FILL_5_NAND2X1_68 ( );
FILL FILL_6_NAND2X1_68 ( );
FILL FILL_0_AND2X2_29 ( );
FILL FILL_1_AND2X2_29 ( );
FILL FILL_2_AND2X2_29 ( );
FILL FILL_3_AND2X2_29 ( );
FILL FILL_4_AND2X2_29 ( );
FILL FILL_5_AND2X2_29 ( );
FILL FILL_6_AND2X2_29 ( );
FILL FILL_7_AND2X2_29 ( );
FILL FILL_8_AND2X2_29 ( );
FILL FILL_0_BUFX2_59 ( );
FILL FILL_1_BUFX2_59 ( );
FILL FILL_2_BUFX2_59 ( );
FILL FILL_3_BUFX2_59 ( );
FILL FILL_4_BUFX2_59 ( );
FILL FILL_5_BUFX2_59 ( );
FILL FILL_6_BUFX2_59 ( );
FILL FILL_0_BUFX2_57 ( );
FILL FILL_1_BUFX2_57 ( );
FILL FILL_2_BUFX2_57 ( );
FILL FILL_3_BUFX2_57 ( );
FILL FILL_4_BUFX2_57 ( );
FILL FILL_5_BUFX2_57 ( );
FILL FILL_6_BUFX2_57 ( );
FILL FILL_0_DFFPOSX1_26 ( );
FILL FILL_1_DFFPOSX1_26 ( );
FILL FILL_2_DFFPOSX1_26 ( );
FILL FILL_3_DFFPOSX1_26 ( );
FILL FILL_4_DFFPOSX1_26 ( );
FILL FILL_5_DFFPOSX1_26 ( );
FILL FILL_6_DFFPOSX1_26 ( );
FILL FILL_7_DFFPOSX1_26 ( );
FILL FILL_8_DFFPOSX1_26 ( );
FILL FILL_9_DFFPOSX1_26 ( );
FILL FILL_10_DFFPOSX1_26 ( );
FILL FILL_11_DFFPOSX1_26 ( );
FILL FILL_12_DFFPOSX1_26 ( );
FILL FILL_13_DFFPOSX1_26 ( );
FILL FILL_14_DFFPOSX1_26 ( );
FILL FILL_15_DFFPOSX1_26 ( );
FILL FILL_16_DFFPOSX1_26 ( );
FILL FILL_17_DFFPOSX1_26 ( );
FILL FILL_18_DFFPOSX1_26 ( );
FILL FILL_19_DFFPOSX1_26 ( );
FILL FILL_20_DFFPOSX1_26 ( );
FILL FILL_21_DFFPOSX1_26 ( );
FILL FILL_22_DFFPOSX1_26 ( );
FILL FILL_23_DFFPOSX1_26 ( );
FILL FILL_24_DFFPOSX1_26 ( );
FILL FILL_25_DFFPOSX1_26 ( );
FILL FILL_26_DFFPOSX1_26 ( );
FILL FILL_27_DFFPOSX1_26 ( );
FILL FILL_0_DFFPOSX1_12 ( );
FILL FILL_1_DFFPOSX1_12 ( );
FILL FILL_2_DFFPOSX1_12 ( );
FILL FILL_3_DFFPOSX1_12 ( );
FILL FILL_4_DFFPOSX1_12 ( );
FILL FILL_5_DFFPOSX1_12 ( );
FILL FILL_6_DFFPOSX1_12 ( );
FILL FILL_7_DFFPOSX1_12 ( );
FILL FILL_8_DFFPOSX1_12 ( );
FILL FILL_9_DFFPOSX1_12 ( );
FILL FILL_10_DFFPOSX1_12 ( );
FILL FILL_11_DFFPOSX1_12 ( );
FILL FILL_12_DFFPOSX1_12 ( );
FILL FILL_13_DFFPOSX1_12 ( );
FILL FILL_14_DFFPOSX1_12 ( );
FILL FILL_15_DFFPOSX1_12 ( );
FILL FILL_16_DFFPOSX1_12 ( );
FILL FILL_17_DFFPOSX1_12 ( );
FILL FILL_18_DFFPOSX1_12 ( );
FILL FILL_19_DFFPOSX1_12 ( );
FILL FILL_20_DFFPOSX1_12 ( );
FILL FILL_21_DFFPOSX1_12 ( );
FILL FILL_22_DFFPOSX1_12 ( );
FILL FILL_23_DFFPOSX1_12 ( );
FILL FILL_24_DFFPOSX1_12 ( );
FILL FILL_25_DFFPOSX1_12 ( );
FILL FILL_26_DFFPOSX1_12 ( );
FILL FILL_27_DFFPOSX1_12 ( );
FILL FILL_0_INVX1_129 ( );
FILL FILL_1_INVX1_129 ( );
FILL FILL_2_INVX1_129 ( );
FILL FILL_3_INVX1_129 ( );
FILL FILL_0_CLKBUF1_43 ( );
FILL FILL_1_CLKBUF1_43 ( );
FILL FILL_2_CLKBUF1_43 ( );
FILL FILL_3_CLKBUF1_43 ( );
FILL FILL_4_CLKBUF1_43 ( );
FILL FILL_5_CLKBUF1_43 ( );
FILL FILL_6_CLKBUF1_43 ( );
FILL FILL_7_CLKBUF1_43 ( );
FILL FILL_8_CLKBUF1_43 ( );
FILL FILL_9_CLKBUF1_43 ( );
FILL FILL_10_CLKBUF1_43 ( );
FILL FILL_11_CLKBUF1_43 ( );
FILL FILL_12_CLKBUF1_43 ( );
FILL FILL_13_CLKBUF1_43 ( );
FILL FILL_14_CLKBUF1_43 ( );
FILL FILL_15_CLKBUF1_43 ( );
FILL FILL_16_CLKBUF1_43 ( );
FILL FILL_17_CLKBUF1_43 ( );
FILL FILL_18_CLKBUF1_43 ( );
FILL FILL_19_CLKBUF1_43 ( );
FILL FILL_20_CLKBUF1_43 ( );
FILL FILL_0_DFFPOSX1_6 ( );
FILL FILL_1_DFFPOSX1_6 ( );
FILL FILL_2_DFFPOSX1_6 ( );
FILL FILL_3_DFFPOSX1_6 ( );
FILL FILL_4_DFFPOSX1_6 ( );
FILL FILL_5_DFFPOSX1_6 ( );
FILL FILL_6_DFFPOSX1_6 ( );
FILL FILL_7_DFFPOSX1_6 ( );
FILL FILL_8_DFFPOSX1_6 ( );
FILL FILL_9_DFFPOSX1_6 ( );
FILL FILL_10_DFFPOSX1_6 ( );
FILL FILL_11_DFFPOSX1_6 ( );
FILL FILL_12_DFFPOSX1_6 ( );
FILL FILL_13_DFFPOSX1_6 ( );
FILL FILL_14_DFFPOSX1_6 ( );
FILL FILL_15_DFFPOSX1_6 ( );
FILL FILL_16_DFFPOSX1_6 ( );
FILL FILL_17_DFFPOSX1_6 ( );
FILL FILL_18_DFFPOSX1_6 ( );
FILL FILL_19_DFFPOSX1_6 ( );
FILL FILL_20_DFFPOSX1_6 ( );
FILL FILL_21_DFFPOSX1_6 ( );
FILL FILL_22_DFFPOSX1_6 ( );
FILL FILL_23_DFFPOSX1_6 ( );
FILL FILL_24_DFFPOSX1_6 ( );
FILL FILL_25_DFFPOSX1_6 ( );
FILL FILL_26_DFFPOSX1_6 ( );
FILL FILL_27_DFFPOSX1_6 ( );
FILL FILL_0_INVX1_38 ( );
FILL FILL_1_INVX1_38 ( );
FILL FILL_2_INVX1_38 ( );
FILL FILL_3_INVX1_38 ( );
FILL FILL_4_INVX1_38 ( );
FILL FILL_0_BUFX2_43 ( );
FILL FILL_1_BUFX2_43 ( );
FILL FILL_2_BUFX2_43 ( );
FILL FILL_3_BUFX2_43 ( );
FILL FILL_4_BUFX2_43 ( );
FILL FILL_5_BUFX2_43 ( );
FILL FILL_6_BUFX2_43 ( );
FILL FILL_0_DFFSR_23 ( );
FILL FILL_1_DFFSR_23 ( );
FILL FILL_2_DFFSR_23 ( );
FILL FILL_3_DFFSR_23 ( );
FILL FILL_4_DFFSR_23 ( );
FILL FILL_5_DFFSR_23 ( );
FILL FILL_6_DFFSR_23 ( );
FILL FILL_7_DFFSR_23 ( );
FILL FILL_8_DFFSR_23 ( );
FILL FILL_9_DFFSR_23 ( );
FILL FILL_10_DFFSR_23 ( );
FILL FILL_11_DFFSR_23 ( );
FILL FILL_12_DFFSR_23 ( );
FILL FILL_13_DFFSR_23 ( );
FILL FILL_14_DFFSR_23 ( );
FILL FILL_15_DFFSR_23 ( );
FILL FILL_16_DFFSR_23 ( );
FILL FILL_17_DFFSR_23 ( );
FILL FILL_18_DFFSR_23 ( );
FILL FILL_19_DFFSR_23 ( );
FILL FILL_20_DFFSR_23 ( );
FILL FILL_21_DFFSR_23 ( );
FILL FILL_22_DFFSR_23 ( );
FILL FILL_23_DFFSR_23 ( );
FILL FILL_24_DFFSR_23 ( );
FILL FILL_25_DFFSR_23 ( );
FILL FILL_26_DFFSR_23 ( );
FILL FILL_27_DFFSR_23 ( );
FILL FILL_28_DFFSR_23 ( );
FILL FILL_29_DFFSR_23 ( );
FILL FILL_30_DFFSR_23 ( );
FILL FILL_31_DFFSR_23 ( );
FILL FILL_32_DFFSR_23 ( );
FILL FILL_33_DFFSR_23 ( );
FILL FILL_34_DFFSR_23 ( );
FILL FILL_35_DFFSR_23 ( );
FILL FILL_36_DFFSR_23 ( );
FILL FILL_37_DFFSR_23 ( );
FILL FILL_38_DFFSR_23 ( );
FILL FILL_39_DFFSR_23 ( );
FILL FILL_40_DFFSR_23 ( );
FILL FILL_41_DFFSR_23 ( );
FILL FILL_42_DFFSR_23 ( );
FILL FILL_43_DFFSR_23 ( );
FILL FILL_44_DFFSR_23 ( );
FILL FILL_45_DFFSR_23 ( );
FILL FILL_46_DFFSR_23 ( );
FILL FILL_47_DFFSR_23 ( );
FILL FILL_48_DFFSR_23 ( );
FILL FILL_49_DFFSR_23 ( );
FILL FILL_50_DFFSR_23 ( );
FILL FILL_0_OAI21X1_20 ( );
FILL FILL_1_OAI21X1_20 ( );
FILL FILL_2_OAI21X1_20 ( );
FILL FILL_3_OAI21X1_20 ( );
FILL FILL_4_OAI21X1_20 ( );
FILL FILL_5_OAI21X1_20 ( );
FILL FILL_6_OAI21X1_20 ( );
FILL FILL_7_OAI21X1_20 ( );
FILL FILL_8_OAI21X1_20 ( );
FILL FILL_9_OAI21X1_20 ( );
FILL FILL_0_NAND3X1_132 ( );
FILL FILL_1_NAND3X1_132 ( );
FILL FILL_2_NAND3X1_132 ( );
FILL FILL_3_NAND3X1_132 ( );
FILL FILL_4_NAND3X1_132 ( );
FILL FILL_5_NAND3X1_132 ( );
FILL FILL_6_NAND3X1_132 ( );
FILL FILL_7_NAND3X1_132 ( );
FILL FILL_8_NAND3X1_132 ( );
FILL FILL_0_DFFSR_252 ( );
FILL FILL_1_DFFSR_252 ( );
FILL FILL_2_DFFSR_252 ( );
FILL FILL_3_DFFSR_252 ( );
FILL FILL_4_DFFSR_252 ( );
FILL FILL_5_DFFSR_252 ( );
FILL FILL_6_DFFSR_252 ( );
FILL FILL_7_DFFSR_252 ( );
FILL FILL_8_DFFSR_252 ( );
FILL FILL_9_DFFSR_252 ( );
FILL FILL_10_DFFSR_252 ( );
FILL FILL_11_DFFSR_252 ( );
FILL FILL_12_DFFSR_252 ( );
FILL FILL_13_DFFSR_252 ( );
FILL FILL_14_DFFSR_252 ( );
FILL FILL_15_DFFSR_252 ( );
FILL FILL_16_DFFSR_252 ( );
FILL FILL_17_DFFSR_252 ( );
FILL FILL_18_DFFSR_252 ( );
FILL FILL_19_DFFSR_252 ( );
FILL FILL_20_DFFSR_252 ( );
FILL FILL_21_DFFSR_252 ( );
FILL FILL_22_DFFSR_252 ( );
FILL FILL_23_DFFSR_252 ( );
FILL FILL_24_DFFSR_252 ( );
FILL FILL_25_DFFSR_252 ( );
FILL FILL_26_DFFSR_252 ( );
FILL FILL_27_DFFSR_252 ( );
FILL FILL_28_DFFSR_252 ( );
FILL FILL_29_DFFSR_252 ( );
FILL FILL_30_DFFSR_252 ( );
FILL FILL_31_DFFSR_252 ( );
FILL FILL_32_DFFSR_252 ( );
FILL FILL_33_DFFSR_252 ( );
FILL FILL_34_DFFSR_252 ( );
FILL FILL_35_DFFSR_252 ( );
FILL FILL_36_DFFSR_252 ( );
FILL FILL_37_DFFSR_252 ( );
FILL FILL_38_DFFSR_252 ( );
FILL FILL_39_DFFSR_252 ( );
FILL FILL_40_DFFSR_252 ( );
FILL FILL_41_DFFSR_252 ( );
FILL FILL_42_DFFSR_252 ( );
FILL FILL_43_DFFSR_252 ( );
FILL FILL_44_DFFSR_252 ( );
FILL FILL_45_DFFSR_252 ( );
FILL FILL_46_DFFSR_252 ( );
FILL FILL_47_DFFSR_252 ( );
FILL FILL_48_DFFSR_252 ( );
FILL FILL_49_DFFSR_252 ( );
FILL FILL_50_DFFSR_252 ( );
FILL FILL_0_NAND2X1_27 ( );
FILL FILL_1_NAND2X1_27 ( );
FILL FILL_2_NAND2X1_27 ( );
FILL FILL_3_NAND2X1_27 ( );
FILL FILL_4_NAND2X1_27 ( );
FILL FILL_5_NAND2X1_27 ( );
FILL FILL_6_NAND2X1_27 ( );
FILL FILL_0_NAND2X1_30 ( );
FILL FILL_1_NAND2X1_30 ( );
FILL FILL_2_NAND2X1_30 ( );
FILL FILL_3_NAND2X1_30 ( );
FILL FILL_4_NAND2X1_30 ( );
FILL FILL_5_NAND2X1_30 ( );
FILL FILL_6_NAND2X1_30 ( );
FILL FILL_0_DFFSR_150 ( );
FILL FILL_1_DFFSR_150 ( );
FILL FILL_2_DFFSR_150 ( );
FILL FILL_3_DFFSR_150 ( );
FILL FILL_4_DFFSR_150 ( );
FILL FILL_5_DFFSR_150 ( );
FILL FILL_6_DFFSR_150 ( );
FILL FILL_7_DFFSR_150 ( );
FILL FILL_8_DFFSR_150 ( );
FILL FILL_9_DFFSR_150 ( );
FILL FILL_10_DFFSR_150 ( );
FILL FILL_11_DFFSR_150 ( );
FILL FILL_12_DFFSR_150 ( );
FILL FILL_13_DFFSR_150 ( );
FILL FILL_14_DFFSR_150 ( );
FILL FILL_15_DFFSR_150 ( );
FILL FILL_16_DFFSR_150 ( );
FILL FILL_17_DFFSR_150 ( );
FILL FILL_18_DFFSR_150 ( );
FILL FILL_19_DFFSR_150 ( );
FILL FILL_20_DFFSR_150 ( );
FILL FILL_21_DFFSR_150 ( );
FILL FILL_22_DFFSR_150 ( );
FILL FILL_23_DFFSR_150 ( );
FILL FILL_24_DFFSR_150 ( );
FILL FILL_25_DFFSR_150 ( );
FILL FILL_26_DFFSR_150 ( );
FILL FILL_27_DFFSR_150 ( );
FILL FILL_28_DFFSR_150 ( );
FILL FILL_29_DFFSR_150 ( );
FILL FILL_30_DFFSR_150 ( );
FILL FILL_31_DFFSR_150 ( );
FILL FILL_32_DFFSR_150 ( );
FILL FILL_33_DFFSR_150 ( );
FILL FILL_34_DFFSR_150 ( );
FILL FILL_35_DFFSR_150 ( );
FILL FILL_36_DFFSR_150 ( );
FILL FILL_37_DFFSR_150 ( );
FILL FILL_38_DFFSR_150 ( );
FILL FILL_39_DFFSR_150 ( );
FILL FILL_40_DFFSR_150 ( );
FILL FILL_41_DFFSR_150 ( );
FILL FILL_42_DFFSR_150 ( );
FILL FILL_43_DFFSR_150 ( );
FILL FILL_44_DFFSR_150 ( );
FILL FILL_45_DFFSR_150 ( );
FILL FILL_46_DFFSR_150 ( );
FILL FILL_47_DFFSR_150 ( );
FILL FILL_48_DFFSR_150 ( );
FILL FILL_49_DFFSR_150 ( );
FILL FILL_50_DFFSR_150 ( );
FILL FILL_0_NAND3X1_103 ( );
FILL FILL_1_NAND3X1_103 ( );
FILL FILL_2_NAND3X1_103 ( );
FILL FILL_3_NAND3X1_103 ( );
FILL FILL_4_NAND3X1_103 ( );
FILL FILL_5_NAND3X1_103 ( );
FILL FILL_6_NAND3X1_103 ( );
FILL FILL_7_NAND3X1_103 ( );
FILL FILL_8_NAND3X1_103 ( );
FILL FILL_9_NAND3X1_103 ( );
FILL FILL_0_NAND3X1_104 ( );
FILL FILL_1_NAND3X1_104 ( );
FILL FILL_2_NAND3X1_104 ( );
FILL FILL_3_NAND3X1_104 ( );
FILL FILL_4_NAND3X1_104 ( );
FILL FILL_5_NAND3X1_104 ( );
FILL FILL_6_NAND3X1_104 ( );
FILL FILL_7_NAND3X1_104 ( );
FILL FILL_8_NAND3X1_104 ( );
FILL FILL_0_NOR2X1_47 ( );
FILL FILL_1_NOR2X1_47 ( );
FILL FILL_2_NOR2X1_47 ( );
FILL FILL_3_NOR2X1_47 ( );
FILL FILL_4_NOR2X1_47 ( );
FILL FILL_5_NOR2X1_47 ( );
FILL FILL_6_NOR2X1_47 ( );
FILL FILL_0_OAI22X1_38 ( );
FILL FILL_1_OAI22X1_38 ( );
FILL FILL_2_OAI22X1_38 ( );
FILL FILL_3_OAI22X1_38 ( );
FILL FILL_4_OAI22X1_38 ( );
FILL FILL_5_OAI22X1_38 ( );
FILL FILL_6_OAI22X1_38 ( );
FILL FILL_7_OAI22X1_38 ( );
FILL FILL_8_OAI22X1_38 ( );
FILL FILL_9_OAI22X1_38 ( );
FILL FILL_10_OAI22X1_38 ( );
FILL FILL_0_INVX1_112 ( );
FILL FILL_1_INVX1_112 ( );
FILL FILL_2_INVX1_112 ( );
FILL FILL_3_INVX1_112 ( );
FILL FILL_4_INVX1_112 ( );
FILL FILL_0_INVX1_91 ( );
FILL FILL_1_INVX1_91 ( );
FILL FILL_2_INVX1_91 ( );
FILL FILL_3_INVX1_91 ( );
FILL FILL_4_INVX1_91 ( );
FILL FILL_0_AOI22X1_13 ( );
FILL FILL_1_AOI22X1_13 ( );
FILL FILL_2_AOI22X1_13 ( );
FILL FILL_3_AOI22X1_13 ( );
FILL FILL_4_AOI22X1_13 ( );
FILL FILL_5_AOI22X1_13 ( );
FILL FILL_6_AOI22X1_13 ( );
FILL FILL_7_AOI22X1_13 ( );
FILL FILL_8_AOI22X1_13 ( );
FILL FILL_9_AOI22X1_13 ( );
FILL FILL_10_AOI22X1_13 ( );
FILL FILL_0_CLKBUF1_12 ( );
FILL FILL_1_CLKBUF1_12 ( );
FILL FILL_2_CLKBUF1_12 ( );
FILL FILL_3_CLKBUF1_12 ( );
FILL FILL_4_CLKBUF1_12 ( );
FILL FILL_5_CLKBUF1_12 ( );
FILL FILL_6_CLKBUF1_12 ( );
FILL FILL_7_CLKBUF1_12 ( );
FILL FILL_8_CLKBUF1_12 ( );
FILL FILL_9_CLKBUF1_12 ( );
FILL FILL_10_CLKBUF1_12 ( );
FILL FILL_11_CLKBUF1_12 ( );
FILL FILL_12_CLKBUF1_12 ( );
FILL FILL_13_CLKBUF1_12 ( );
FILL FILL_14_CLKBUF1_12 ( );
FILL FILL_15_CLKBUF1_12 ( );
FILL FILL_16_CLKBUF1_12 ( );
FILL FILL_17_CLKBUF1_12 ( );
FILL FILL_18_CLKBUF1_12 ( );
FILL FILL_19_CLKBUF1_12 ( );
FILL FILL_20_CLKBUF1_12 ( );
FILL FILL_0_INVX1_92 ( );
FILL FILL_1_INVX1_92 ( );
FILL FILL_2_INVX1_92 ( );
FILL FILL_3_INVX1_92 ( );
FILL FILL_4_INVX1_92 ( );
FILL FILL_0_OAI21X1_72 ( );
FILL FILL_1_OAI21X1_72 ( );
FILL FILL_2_OAI21X1_72 ( );
FILL FILL_3_OAI21X1_72 ( );
FILL FILL_4_OAI21X1_72 ( );
FILL FILL_5_OAI21X1_72 ( );
FILL FILL_6_OAI21X1_72 ( );
FILL FILL_7_OAI21X1_72 ( );
FILL FILL_8_OAI21X1_72 ( );
FILL FILL_0_OAI21X1_69 ( );
FILL FILL_1_OAI21X1_69 ( );
FILL FILL_2_OAI21X1_69 ( );
FILL FILL_3_OAI21X1_69 ( );
FILL FILL_4_OAI21X1_69 ( );
FILL FILL_5_OAI21X1_69 ( );
FILL FILL_6_OAI21X1_69 ( );
FILL FILL_7_OAI21X1_69 ( );
FILL FILL_8_OAI21X1_69 ( );
FILL FILL_0_OAI21X1_70 ( );
FILL FILL_1_OAI21X1_70 ( );
FILL FILL_2_OAI21X1_70 ( );
FILL FILL_3_OAI21X1_70 ( );
FILL FILL_4_OAI21X1_70 ( );
FILL FILL_5_OAI21X1_70 ( );
FILL FILL_6_OAI21X1_70 ( );
FILL FILL_7_OAI21X1_70 ( );
FILL FILL_8_OAI21X1_70 ( );
FILL FILL_0_OAI22X1_50 ( );
FILL FILL_1_OAI22X1_50 ( );
FILL FILL_2_OAI22X1_50 ( );
FILL FILL_3_OAI22X1_50 ( );
FILL FILL_4_OAI22X1_50 ( );
FILL FILL_5_OAI22X1_50 ( );
FILL FILL_6_OAI22X1_50 ( );
FILL FILL_7_OAI22X1_50 ( );
FILL FILL_8_OAI22X1_50 ( );
FILL FILL_9_OAI22X1_50 ( );
FILL FILL_10_OAI22X1_50 ( );
FILL FILL_0_NAND2X1_69 ( );
FILL FILL_1_NAND2X1_69 ( );
FILL FILL_2_NAND2X1_69 ( );
FILL FILL_3_NAND2X1_69 ( );
FILL FILL_4_NAND2X1_69 ( );
FILL FILL_5_NAND2X1_69 ( );
FILL FILL_6_NAND2X1_69 ( );
FILL FILL_0_NAND3X1_157 ( );
FILL FILL_1_NAND3X1_157 ( );
FILL FILL_2_NAND3X1_157 ( );
FILL FILL_3_NAND3X1_157 ( );
FILL FILL_4_NAND3X1_157 ( );
FILL FILL_5_NAND3X1_157 ( );
FILL FILL_6_NAND3X1_157 ( );
FILL FILL_7_NAND3X1_157 ( );
FILL FILL_8_NAND3X1_157 ( );
FILL FILL_0_NAND2X1_76 ( );
FILL FILL_1_NAND2X1_76 ( );
FILL FILL_2_NAND2X1_76 ( );
FILL FILL_3_NAND2X1_76 ( );
FILL FILL_4_NAND2X1_76 ( );
FILL FILL_5_NAND2X1_76 ( );
FILL FILL_6_NAND2X1_76 ( );
FILL FILL_0_DFFSR_272 ( );
FILL FILL_1_DFFSR_272 ( );
FILL FILL_2_DFFSR_272 ( );
FILL FILL_3_DFFSR_272 ( );
FILL FILL_4_DFFSR_272 ( );
FILL FILL_5_DFFSR_272 ( );
FILL FILL_6_DFFSR_272 ( );
FILL FILL_7_DFFSR_272 ( );
FILL FILL_8_DFFSR_272 ( );
FILL FILL_9_DFFSR_272 ( );
FILL FILL_10_DFFSR_272 ( );
FILL FILL_11_DFFSR_272 ( );
FILL FILL_12_DFFSR_272 ( );
FILL FILL_13_DFFSR_272 ( );
FILL FILL_14_DFFSR_272 ( );
FILL FILL_15_DFFSR_272 ( );
FILL FILL_16_DFFSR_272 ( );
FILL FILL_17_DFFSR_272 ( );
FILL FILL_18_DFFSR_272 ( );
FILL FILL_19_DFFSR_272 ( );
FILL FILL_20_DFFSR_272 ( );
FILL FILL_21_DFFSR_272 ( );
FILL FILL_22_DFFSR_272 ( );
FILL FILL_23_DFFSR_272 ( );
FILL FILL_24_DFFSR_272 ( );
FILL FILL_25_DFFSR_272 ( );
FILL FILL_26_DFFSR_272 ( );
FILL FILL_27_DFFSR_272 ( );
FILL FILL_28_DFFSR_272 ( );
FILL FILL_29_DFFSR_272 ( );
FILL FILL_30_DFFSR_272 ( );
FILL FILL_31_DFFSR_272 ( );
FILL FILL_32_DFFSR_272 ( );
FILL FILL_33_DFFSR_272 ( );
FILL FILL_34_DFFSR_272 ( );
FILL FILL_35_DFFSR_272 ( );
FILL FILL_36_DFFSR_272 ( );
FILL FILL_37_DFFSR_272 ( );
FILL FILL_38_DFFSR_272 ( );
FILL FILL_39_DFFSR_272 ( );
FILL FILL_40_DFFSR_272 ( );
FILL FILL_41_DFFSR_272 ( );
FILL FILL_42_DFFSR_272 ( );
FILL FILL_43_DFFSR_272 ( );
FILL FILL_44_DFFSR_272 ( );
FILL FILL_45_DFFSR_272 ( );
FILL FILL_46_DFFSR_272 ( );
FILL FILL_47_DFFSR_272 ( );
FILL FILL_48_DFFSR_272 ( );
FILL FILL_49_DFFSR_272 ( );
FILL FILL_50_DFFSR_272 ( );
FILL FILL_0_AOI21X1_62 ( );
FILL FILL_1_AOI21X1_62 ( );
FILL FILL_2_AOI21X1_62 ( );
FILL FILL_3_AOI21X1_62 ( );
FILL FILL_4_AOI21X1_62 ( );
FILL FILL_5_AOI21X1_62 ( );
FILL FILL_6_AOI21X1_62 ( );
FILL FILL_7_AOI21X1_62 ( );
FILL FILL_8_AOI21X1_62 ( );
FILL FILL_9_AOI21X1_62 ( );
FILL FILL_0_AOI21X1_5 ( );
FILL FILL_1_AOI21X1_5 ( );
FILL FILL_2_AOI21X1_5 ( );
FILL FILL_3_AOI21X1_5 ( );
FILL FILL_4_AOI21X1_5 ( );
FILL FILL_5_AOI21X1_5 ( );
FILL FILL_6_AOI21X1_5 ( );
FILL FILL_7_AOI21X1_5 ( );
FILL FILL_8_AOI21X1_5 ( );
FILL FILL_0_XOR2X1_12 ( );
FILL FILL_1_XOR2X1_12 ( );
FILL FILL_2_XOR2X1_12 ( );
FILL FILL_3_XOR2X1_12 ( );
FILL FILL_4_XOR2X1_12 ( );
FILL FILL_5_XOR2X1_12 ( );
FILL FILL_6_XOR2X1_12 ( );
FILL FILL_7_XOR2X1_12 ( );
FILL FILL_8_XOR2X1_12 ( );
FILL FILL_9_XOR2X1_12 ( );
FILL FILL_10_XOR2X1_12 ( );
FILL FILL_11_XOR2X1_12 ( );
FILL FILL_12_XOR2X1_12 ( );
FILL FILL_13_XOR2X1_12 ( );
FILL FILL_14_XOR2X1_12 ( );
FILL FILL_15_XOR2X1_12 ( );
FILL FILL_0_NOR2X1_63 ( );
FILL FILL_1_NOR2X1_63 ( );
FILL FILL_2_NOR2X1_63 ( );
FILL FILL_3_NOR2X1_63 ( );
FILL FILL_4_NOR2X1_63 ( );
FILL FILL_5_NOR2X1_63 ( );
FILL FILL_6_NOR2X1_63 ( );
FILL FILL_0_AOI21X1_65 ( );
FILL FILL_1_AOI21X1_65 ( );
FILL FILL_2_AOI21X1_65 ( );
FILL FILL_3_AOI21X1_65 ( );
FILL FILL_4_AOI21X1_65 ( );
FILL FILL_5_AOI21X1_65 ( );
FILL FILL_6_AOI21X1_65 ( );
FILL FILL_7_AOI21X1_65 ( );
FILL FILL_8_AOI21X1_65 ( );
FILL FILL_0_DFFSR_116 ( );
FILL FILL_1_DFFSR_116 ( );
FILL FILL_2_DFFSR_116 ( );
FILL FILL_3_DFFSR_116 ( );
FILL FILL_4_DFFSR_116 ( );
FILL FILL_5_DFFSR_116 ( );
FILL FILL_6_DFFSR_116 ( );
FILL FILL_7_DFFSR_116 ( );
FILL FILL_8_DFFSR_116 ( );
FILL FILL_9_DFFSR_116 ( );
FILL FILL_10_DFFSR_116 ( );
FILL FILL_11_DFFSR_116 ( );
FILL FILL_12_DFFSR_116 ( );
FILL FILL_13_DFFSR_116 ( );
FILL FILL_14_DFFSR_116 ( );
FILL FILL_15_DFFSR_116 ( );
FILL FILL_16_DFFSR_116 ( );
FILL FILL_17_DFFSR_116 ( );
FILL FILL_18_DFFSR_116 ( );
FILL FILL_19_DFFSR_116 ( );
FILL FILL_20_DFFSR_116 ( );
FILL FILL_21_DFFSR_116 ( );
FILL FILL_22_DFFSR_116 ( );
FILL FILL_23_DFFSR_116 ( );
FILL FILL_24_DFFSR_116 ( );
FILL FILL_25_DFFSR_116 ( );
FILL FILL_26_DFFSR_116 ( );
FILL FILL_27_DFFSR_116 ( );
FILL FILL_28_DFFSR_116 ( );
FILL FILL_29_DFFSR_116 ( );
FILL FILL_30_DFFSR_116 ( );
FILL FILL_31_DFFSR_116 ( );
FILL FILL_32_DFFSR_116 ( );
FILL FILL_33_DFFSR_116 ( );
FILL FILL_34_DFFSR_116 ( );
FILL FILL_35_DFFSR_116 ( );
FILL FILL_36_DFFSR_116 ( );
FILL FILL_37_DFFSR_116 ( );
FILL FILL_38_DFFSR_116 ( );
FILL FILL_39_DFFSR_116 ( );
FILL FILL_40_DFFSR_116 ( );
FILL FILL_41_DFFSR_116 ( );
FILL FILL_42_DFFSR_116 ( );
FILL FILL_43_DFFSR_116 ( );
FILL FILL_44_DFFSR_116 ( );
FILL FILL_45_DFFSR_116 ( );
FILL FILL_46_DFFSR_116 ( );
FILL FILL_47_DFFSR_116 ( );
FILL FILL_48_DFFSR_116 ( );
FILL FILL_49_DFFSR_116 ( );
FILL FILL_50_DFFSR_116 ( );
FILL FILL_0_BUFX2_88 ( );
FILL FILL_1_BUFX2_88 ( );
FILL FILL_2_BUFX2_88 ( );
FILL FILL_3_BUFX2_88 ( );
FILL FILL_4_BUFX2_88 ( );
FILL FILL_5_BUFX2_88 ( );
FILL FILL_6_BUFX2_88 ( );
FILL FILL_0_AND2X2_42 ( );
FILL FILL_1_AND2X2_42 ( );
FILL FILL_2_AND2X2_42 ( );
FILL FILL_3_AND2X2_42 ( );
FILL FILL_4_AND2X2_42 ( );
FILL FILL_5_AND2X2_42 ( );
FILL FILL_6_AND2X2_42 ( );
FILL FILL_7_AND2X2_42 ( );
FILL FILL_8_AND2X2_42 ( );
FILL FILL_9_AND2X2_42 ( );
FILL FILL_0_DFFSR_120 ( );
FILL FILL_1_DFFSR_120 ( );
FILL FILL_2_DFFSR_120 ( );
FILL FILL_3_DFFSR_120 ( );
FILL FILL_4_DFFSR_120 ( );
FILL FILL_5_DFFSR_120 ( );
FILL FILL_6_DFFSR_120 ( );
FILL FILL_7_DFFSR_120 ( );
FILL FILL_8_DFFSR_120 ( );
FILL FILL_9_DFFSR_120 ( );
FILL FILL_10_DFFSR_120 ( );
FILL FILL_11_DFFSR_120 ( );
FILL FILL_12_DFFSR_120 ( );
FILL FILL_13_DFFSR_120 ( );
FILL FILL_14_DFFSR_120 ( );
FILL FILL_15_DFFSR_120 ( );
FILL FILL_16_DFFSR_120 ( );
FILL FILL_17_DFFSR_120 ( );
FILL FILL_18_DFFSR_120 ( );
FILL FILL_19_DFFSR_120 ( );
FILL FILL_20_DFFSR_120 ( );
FILL FILL_21_DFFSR_120 ( );
FILL FILL_22_DFFSR_120 ( );
FILL FILL_23_DFFSR_120 ( );
FILL FILL_24_DFFSR_120 ( );
FILL FILL_25_DFFSR_120 ( );
FILL FILL_26_DFFSR_120 ( );
FILL FILL_27_DFFSR_120 ( );
FILL FILL_28_DFFSR_120 ( );
FILL FILL_29_DFFSR_120 ( );
FILL FILL_30_DFFSR_120 ( );
FILL FILL_31_DFFSR_120 ( );
FILL FILL_32_DFFSR_120 ( );
FILL FILL_33_DFFSR_120 ( );
FILL FILL_34_DFFSR_120 ( );
FILL FILL_35_DFFSR_120 ( );
FILL FILL_36_DFFSR_120 ( );
FILL FILL_37_DFFSR_120 ( );
FILL FILL_38_DFFSR_120 ( );
FILL FILL_39_DFFSR_120 ( );
FILL FILL_40_DFFSR_120 ( );
FILL FILL_41_DFFSR_120 ( );
FILL FILL_42_DFFSR_120 ( );
FILL FILL_43_DFFSR_120 ( );
FILL FILL_44_DFFSR_120 ( );
FILL FILL_45_DFFSR_120 ( );
FILL FILL_46_DFFSR_120 ( );
FILL FILL_47_DFFSR_120 ( );
FILL FILL_48_DFFSR_120 ( );
FILL FILL_49_DFFSR_120 ( );
FILL FILL_50_DFFSR_120 ( );
FILL FILL_51_DFFSR_120 ( );
FILL FILL_0_INVX1_126 ( );
FILL FILL_1_INVX1_126 ( );
FILL FILL_2_INVX1_126 ( );
FILL FILL_3_INVX1_126 ( );
FILL FILL_0_AND2X2_15 ( );
FILL FILL_1_AND2X2_15 ( );
FILL FILL_2_AND2X2_15 ( );
FILL FILL_3_AND2X2_15 ( );
FILL FILL_4_AND2X2_15 ( );
FILL FILL_5_AND2X2_15 ( );
FILL FILL_6_AND2X2_15 ( );
FILL FILL_7_AND2X2_15 ( );
FILL FILL_8_AND2X2_15 ( );
FILL FILL_9_AND2X2_15 ( );
FILL FILL_0_NOR2X1_30 ( );
FILL FILL_1_NOR2X1_30 ( );
FILL FILL_2_NOR2X1_30 ( );
FILL FILL_3_NOR2X1_30 ( );
FILL FILL_4_NOR2X1_30 ( );
FILL FILL_5_NOR2X1_30 ( );
FILL FILL_6_NOR2X1_30 ( );
FILL FILL_0_NOR2X1_33 ( );
FILL FILL_1_NOR2X1_33 ( );
FILL FILL_2_NOR2X1_33 ( );
FILL FILL_3_NOR2X1_33 ( );
FILL FILL_4_NOR2X1_33 ( );
FILL FILL_5_NOR2X1_33 ( );
FILL FILL_6_NOR2X1_33 ( );
FILL FILL_0_NAND2X1_29 ( );
FILL FILL_1_NAND2X1_29 ( );
FILL FILL_2_NAND2X1_29 ( );
FILL FILL_3_NAND2X1_29 ( );
FILL FILL_4_NAND2X1_29 ( );
FILL FILL_5_NAND2X1_29 ( );
FILL FILL_6_NAND2X1_29 ( );
FILL FILL_0_NAND2X1_31 ( );
FILL FILL_1_NAND2X1_31 ( );
FILL FILL_2_NAND2X1_31 ( );
FILL FILL_3_NAND2X1_31 ( );
FILL FILL_4_NAND2X1_31 ( );
FILL FILL_5_NAND2X1_31 ( );
FILL FILL_6_NAND2X1_31 ( );
FILL FILL_0_NAND3X1_106 ( );
FILL FILL_1_NAND3X1_106 ( );
FILL FILL_2_NAND3X1_106 ( );
FILL FILL_3_NAND3X1_106 ( );
FILL FILL_4_NAND3X1_106 ( );
FILL FILL_5_NAND3X1_106 ( );
FILL FILL_6_NAND3X1_106 ( );
FILL FILL_7_NAND3X1_106 ( );
FILL FILL_8_NAND3X1_106 ( );
FILL FILL_9_NAND3X1_106 ( );
FILL FILL_0_DFFSR_158 ( );
FILL FILL_1_DFFSR_158 ( );
FILL FILL_2_DFFSR_158 ( );
FILL FILL_3_DFFSR_158 ( );
FILL FILL_4_DFFSR_158 ( );
FILL FILL_5_DFFSR_158 ( );
FILL FILL_6_DFFSR_158 ( );
FILL FILL_7_DFFSR_158 ( );
FILL FILL_8_DFFSR_158 ( );
FILL FILL_9_DFFSR_158 ( );
FILL FILL_10_DFFSR_158 ( );
FILL FILL_11_DFFSR_158 ( );
FILL FILL_12_DFFSR_158 ( );
FILL FILL_13_DFFSR_158 ( );
FILL FILL_14_DFFSR_158 ( );
FILL FILL_15_DFFSR_158 ( );
FILL FILL_16_DFFSR_158 ( );
FILL FILL_17_DFFSR_158 ( );
FILL FILL_18_DFFSR_158 ( );
FILL FILL_19_DFFSR_158 ( );
FILL FILL_20_DFFSR_158 ( );
FILL FILL_21_DFFSR_158 ( );
FILL FILL_22_DFFSR_158 ( );
FILL FILL_23_DFFSR_158 ( );
FILL FILL_24_DFFSR_158 ( );
FILL FILL_25_DFFSR_158 ( );
FILL FILL_26_DFFSR_158 ( );
FILL FILL_27_DFFSR_158 ( );
FILL FILL_28_DFFSR_158 ( );
FILL FILL_29_DFFSR_158 ( );
FILL FILL_30_DFFSR_158 ( );
FILL FILL_31_DFFSR_158 ( );
FILL FILL_32_DFFSR_158 ( );
FILL FILL_33_DFFSR_158 ( );
FILL FILL_34_DFFSR_158 ( );
FILL FILL_35_DFFSR_158 ( );
FILL FILL_36_DFFSR_158 ( );
FILL FILL_37_DFFSR_158 ( );
FILL FILL_38_DFFSR_158 ( );
FILL FILL_39_DFFSR_158 ( );
FILL FILL_40_DFFSR_158 ( );
FILL FILL_41_DFFSR_158 ( );
FILL FILL_42_DFFSR_158 ( );
FILL FILL_43_DFFSR_158 ( );
FILL FILL_44_DFFSR_158 ( );
FILL FILL_45_DFFSR_158 ( );
FILL FILL_46_DFFSR_158 ( );
FILL FILL_47_DFFSR_158 ( );
FILL FILL_48_DFFSR_158 ( );
FILL FILL_49_DFFSR_158 ( );
FILL FILL_50_DFFSR_158 ( );
FILL FILL_51_DFFSR_158 ( );
FILL FILL_0_NAND3X1_102 ( );
FILL FILL_1_NAND3X1_102 ( );
FILL FILL_2_NAND3X1_102 ( );
FILL FILL_3_NAND3X1_102 ( );
FILL FILL_4_NAND3X1_102 ( );
FILL FILL_5_NAND3X1_102 ( );
FILL FILL_6_NAND3X1_102 ( );
FILL FILL_7_NAND3X1_102 ( );
FILL FILL_8_NAND3X1_102 ( );
FILL FILL_9_NAND3X1_102 ( );
FILL FILL_0_OAI22X1_28 ( );
FILL FILL_1_OAI22X1_28 ( );
FILL FILL_2_OAI22X1_28 ( );
FILL FILL_3_OAI22X1_28 ( );
FILL FILL_4_OAI22X1_28 ( );
FILL FILL_5_OAI22X1_28 ( );
FILL FILL_6_OAI22X1_28 ( );
FILL FILL_7_OAI22X1_28 ( );
FILL FILL_8_OAI22X1_28 ( );
FILL FILL_9_OAI22X1_28 ( );
FILL FILL_10_OAI22X1_28 ( );
FILL FILL_0_INVX1_69 ( );
FILL FILL_1_INVX1_69 ( );
FILL FILL_2_INVX1_69 ( );
FILL FILL_3_INVX1_69 ( );
FILL FILL_4_INVX1_69 ( );
FILL FILL_0_OAI22X1_37 ( );
FILL FILL_1_OAI22X1_37 ( );
FILL FILL_2_OAI22X1_37 ( );
FILL FILL_3_OAI22X1_37 ( );
FILL FILL_4_OAI22X1_37 ( );
FILL FILL_5_OAI22X1_37 ( );
FILL FILL_6_OAI22X1_37 ( );
FILL FILL_7_OAI22X1_37 ( );
FILL FILL_8_OAI22X1_37 ( );
FILL FILL_9_OAI22X1_37 ( );
FILL FILL_10_OAI22X1_37 ( );
FILL FILL_0_INVX1_93 ( );
FILL FILL_1_INVX1_93 ( );
FILL FILL_2_INVX1_93 ( );
FILL FILL_3_INVX1_93 ( );
FILL FILL_4_INVX1_93 ( );
FILL FILL_0_DFFSR_213 ( );
FILL FILL_1_DFFSR_213 ( );
FILL FILL_2_DFFSR_213 ( );
FILL FILL_3_DFFSR_213 ( );
FILL FILL_4_DFFSR_213 ( );
FILL FILL_5_DFFSR_213 ( );
FILL FILL_6_DFFSR_213 ( );
FILL FILL_7_DFFSR_213 ( );
FILL FILL_8_DFFSR_213 ( );
FILL FILL_9_DFFSR_213 ( );
FILL FILL_10_DFFSR_213 ( );
FILL FILL_11_DFFSR_213 ( );
FILL FILL_12_DFFSR_213 ( );
FILL FILL_13_DFFSR_213 ( );
FILL FILL_14_DFFSR_213 ( );
FILL FILL_15_DFFSR_213 ( );
FILL FILL_16_DFFSR_213 ( );
FILL FILL_17_DFFSR_213 ( );
FILL FILL_18_DFFSR_213 ( );
FILL FILL_19_DFFSR_213 ( );
FILL FILL_20_DFFSR_213 ( );
FILL FILL_21_DFFSR_213 ( );
FILL FILL_22_DFFSR_213 ( );
FILL FILL_23_DFFSR_213 ( );
FILL FILL_24_DFFSR_213 ( );
FILL FILL_25_DFFSR_213 ( );
FILL FILL_26_DFFSR_213 ( );
FILL FILL_27_DFFSR_213 ( );
FILL FILL_28_DFFSR_213 ( );
FILL FILL_29_DFFSR_213 ( );
FILL FILL_30_DFFSR_213 ( );
FILL FILL_31_DFFSR_213 ( );
FILL FILL_32_DFFSR_213 ( );
FILL FILL_33_DFFSR_213 ( );
FILL FILL_34_DFFSR_213 ( );
FILL FILL_35_DFFSR_213 ( );
FILL FILL_36_DFFSR_213 ( );
FILL FILL_37_DFFSR_213 ( );
FILL FILL_38_DFFSR_213 ( );
FILL FILL_39_DFFSR_213 ( );
FILL FILL_40_DFFSR_213 ( );
FILL FILL_41_DFFSR_213 ( );
FILL FILL_42_DFFSR_213 ( );
FILL FILL_43_DFFSR_213 ( );
FILL FILL_44_DFFSR_213 ( );
FILL FILL_45_DFFSR_213 ( );
FILL FILL_46_DFFSR_213 ( );
FILL FILL_47_DFFSR_213 ( );
FILL FILL_48_DFFSR_213 ( );
FILL FILL_49_DFFSR_213 ( );
FILL FILL_50_DFFSR_213 ( );
FILL FILL_0_INVX1_159 ( );
FILL FILL_1_INVX1_159 ( );
FILL FILL_2_INVX1_159 ( );
FILL FILL_3_INVX1_159 ( );
FILL FILL_4_INVX1_159 ( );
FILL FILL_0_OAI21X1_62 ( );
FILL FILL_1_OAI21X1_62 ( );
FILL FILL_2_OAI21X1_62 ( );
FILL FILL_3_OAI21X1_62 ( );
FILL FILL_4_OAI21X1_62 ( );
FILL FILL_5_OAI21X1_62 ( );
FILL FILL_6_OAI21X1_62 ( );
FILL FILL_7_OAI21X1_62 ( );
FILL FILL_8_OAI21X1_62 ( );
FILL FILL_0_INVX1_134 ( );
FILL FILL_1_INVX1_134 ( );
FILL FILL_2_INVX1_134 ( );
FILL FILL_3_INVX1_134 ( );
FILL FILL_4_INVX1_134 ( );
FILL FILL_0_OAI21X1_71 ( );
FILL FILL_1_OAI21X1_71 ( );
FILL FILL_2_OAI21X1_71 ( );
FILL FILL_3_OAI21X1_71 ( );
FILL FILL_4_OAI21X1_71 ( );
FILL FILL_5_OAI21X1_71 ( );
FILL FILL_6_OAI21X1_71 ( );
FILL FILL_7_OAI21X1_71 ( );
FILL FILL_8_OAI21X1_71 ( );
FILL FILL_9_OAI21X1_71 ( );
FILL FILL_0_AOI22X1_22 ( );
FILL FILL_1_AOI22X1_22 ( );
FILL FILL_2_AOI22X1_22 ( );
FILL FILL_3_AOI22X1_22 ( );
FILL FILL_4_AOI22X1_22 ( );
FILL FILL_5_AOI22X1_22 ( );
FILL FILL_6_AOI22X1_22 ( );
FILL FILL_7_AOI22X1_22 ( );
FILL FILL_8_AOI22X1_22 ( );
FILL FILL_9_AOI22X1_22 ( );
FILL FILL_10_AOI22X1_22 ( );
FILL FILL_11_AOI22X1_22 ( );
FILL FILL_0_INVX1_146 ( );
FILL FILL_1_INVX1_146 ( );
FILL FILL_2_INVX1_146 ( );
FILL FILL_3_INVX1_146 ( );
FILL FILL_0_NAND2X1_75 ( );
FILL FILL_1_NAND2X1_75 ( );
FILL FILL_2_NAND2X1_75 ( );
FILL FILL_3_NAND2X1_75 ( );
FILL FILL_4_NAND2X1_75 ( );
FILL FILL_5_NAND2X1_75 ( );
FILL FILL_6_NAND2X1_75 ( );
FILL FILL_0_OAI21X1_33 ( );
FILL FILL_1_OAI21X1_33 ( );
FILL FILL_2_OAI21X1_33 ( );
FILL FILL_3_OAI21X1_33 ( );
FILL FILL_4_OAI21X1_33 ( );
FILL FILL_5_OAI21X1_33 ( );
FILL FILL_6_OAI21X1_33 ( );
FILL FILL_7_OAI21X1_33 ( );
FILL FILL_8_OAI21X1_33 ( );
FILL FILL_9_OAI21X1_33 ( );
FILL FILL_0_AOI21X1_43 ( );
FILL FILL_1_AOI21X1_43 ( );
FILL FILL_2_AOI21X1_43 ( );
FILL FILL_3_AOI21X1_43 ( );
FILL FILL_4_AOI21X1_43 ( );
FILL FILL_5_AOI21X1_43 ( );
FILL FILL_6_AOI21X1_43 ( );
FILL FILL_7_AOI21X1_43 ( );
FILL FILL_8_AOI21X1_43 ( );
FILL FILL_0_NAND2X1_131 ( );
FILL FILL_1_NAND2X1_131 ( );
FILL FILL_2_NAND2X1_131 ( );
FILL FILL_3_NAND2X1_131 ( );
FILL FILL_4_NAND2X1_131 ( );
FILL FILL_5_NAND2X1_131 ( );
FILL FILL_6_NAND2X1_131 ( );
FILL FILL_0_OAI21X1_100 ( );
FILL FILL_1_OAI21X1_100 ( );
FILL FILL_2_OAI21X1_100 ( );
FILL FILL_3_OAI21X1_100 ( );
FILL FILL_4_OAI21X1_100 ( );
FILL FILL_5_OAI21X1_100 ( );
FILL FILL_6_OAI21X1_100 ( );
FILL FILL_7_OAI21X1_100 ( );
FILL FILL_8_OAI21X1_100 ( );
FILL FILL_9_OAI21X1_100 ( );
FILL FILL_0_INVX1_197 ( );
FILL FILL_1_INVX1_197 ( );
FILL FILL_2_INVX1_197 ( );
FILL FILL_3_INVX1_197 ( );
FILL FILL_0_NOR2X1_76 ( );
FILL FILL_1_NOR2X1_76 ( );
FILL FILL_2_NOR2X1_76 ( );
FILL FILL_3_NOR2X1_76 ( );
FILL FILL_4_NOR2X1_76 ( );
FILL FILL_5_NOR2X1_76 ( );
FILL FILL_6_NOR2X1_76 ( );
FILL FILL_0_CLKBUF1_48 ( );
FILL FILL_1_CLKBUF1_48 ( );
FILL FILL_2_CLKBUF1_48 ( );
FILL FILL_3_CLKBUF1_48 ( );
FILL FILL_4_CLKBUF1_48 ( );
FILL FILL_5_CLKBUF1_48 ( );
FILL FILL_6_CLKBUF1_48 ( );
FILL FILL_7_CLKBUF1_48 ( );
FILL FILL_8_CLKBUF1_48 ( );
FILL FILL_9_CLKBUF1_48 ( );
FILL FILL_10_CLKBUF1_48 ( );
FILL FILL_11_CLKBUF1_48 ( );
FILL FILL_12_CLKBUF1_48 ( );
FILL FILL_13_CLKBUF1_48 ( );
FILL FILL_14_CLKBUF1_48 ( );
FILL FILL_15_CLKBUF1_48 ( );
FILL FILL_16_CLKBUF1_48 ( );
FILL FILL_17_CLKBUF1_48 ( );
FILL FILL_18_CLKBUF1_48 ( );
FILL FILL_19_CLKBUF1_48 ( );
FILL FILL_0_BUFX2_44 ( );
FILL FILL_1_BUFX2_44 ( );
FILL FILL_2_BUFX2_44 ( );
FILL FILL_3_BUFX2_44 ( );
FILL FILL_4_BUFX2_44 ( );
FILL FILL_5_BUFX2_44 ( );
FILL FILL_6_BUFX2_44 ( );
FILL FILL_0_NAND2X1_12 ( );
FILL FILL_1_NAND2X1_12 ( );
FILL FILL_2_NAND2X1_12 ( );
FILL FILL_3_NAND2X1_12 ( );
FILL FILL_4_NAND2X1_12 ( );
FILL FILL_5_NAND2X1_12 ( );
FILL FILL_6_NAND2X1_12 ( );
FILL FILL_0_NOR3X1_1 ( );
FILL FILL_1_NOR3X1_1 ( );
FILL FILL_2_NOR3X1_1 ( );
FILL FILL_3_NOR3X1_1 ( );
FILL FILL_4_NOR3X1_1 ( );
FILL FILL_5_NOR3X1_1 ( );
FILL FILL_6_NOR3X1_1 ( );
FILL FILL_7_NOR3X1_1 ( );
FILL FILL_8_NOR3X1_1 ( );
FILL FILL_9_NOR3X1_1 ( );
FILL FILL_10_NOR3X1_1 ( );
FILL FILL_11_NOR3X1_1 ( );
FILL FILL_12_NOR3X1_1 ( );
FILL FILL_13_NOR3X1_1 ( );
FILL FILL_14_NOR3X1_1 ( );
FILL FILL_15_NOR3X1_1 ( );
FILL FILL_16_NOR3X1_1 ( );
FILL FILL_17_NOR3X1_1 ( );
FILL FILL_18_NOR3X1_1 ( );
FILL FILL_0_INVX1_3 ( );
FILL FILL_1_INVX1_3 ( );
FILL FILL_2_INVX1_3 ( );
FILL FILL_3_INVX1_3 ( );
FILL FILL_0_NAND3X1_248 ( );
FILL FILL_1_NAND3X1_248 ( );
FILL FILL_2_NAND3X1_248 ( );
FILL FILL_3_NAND3X1_248 ( );
FILL FILL_4_NAND3X1_248 ( );
FILL FILL_5_NAND3X1_248 ( );
FILL FILL_6_NAND3X1_248 ( );
FILL FILL_7_NAND3X1_248 ( );
FILL FILL_8_NAND3X1_248 ( );
FILL FILL_9_NAND3X1_248 ( );
FILL FILL_0_DFFSR_39 ( );
FILL FILL_1_DFFSR_39 ( );
FILL FILL_2_DFFSR_39 ( );
FILL FILL_3_DFFSR_39 ( );
FILL FILL_4_DFFSR_39 ( );
FILL FILL_5_DFFSR_39 ( );
FILL FILL_6_DFFSR_39 ( );
FILL FILL_7_DFFSR_39 ( );
FILL FILL_8_DFFSR_39 ( );
FILL FILL_9_DFFSR_39 ( );
FILL FILL_10_DFFSR_39 ( );
FILL FILL_11_DFFSR_39 ( );
FILL FILL_12_DFFSR_39 ( );
FILL FILL_13_DFFSR_39 ( );
FILL FILL_14_DFFSR_39 ( );
FILL FILL_15_DFFSR_39 ( );
FILL FILL_16_DFFSR_39 ( );
FILL FILL_17_DFFSR_39 ( );
FILL FILL_18_DFFSR_39 ( );
FILL FILL_19_DFFSR_39 ( );
FILL FILL_20_DFFSR_39 ( );
FILL FILL_21_DFFSR_39 ( );
FILL FILL_22_DFFSR_39 ( );
FILL FILL_23_DFFSR_39 ( );
FILL FILL_24_DFFSR_39 ( );
FILL FILL_25_DFFSR_39 ( );
FILL FILL_26_DFFSR_39 ( );
FILL FILL_27_DFFSR_39 ( );
FILL FILL_28_DFFSR_39 ( );
FILL FILL_29_DFFSR_39 ( );
FILL FILL_30_DFFSR_39 ( );
FILL FILL_31_DFFSR_39 ( );
FILL FILL_32_DFFSR_39 ( );
FILL FILL_33_DFFSR_39 ( );
FILL FILL_34_DFFSR_39 ( );
FILL FILL_35_DFFSR_39 ( );
FILL FILL_36_DFFSR_39 ( );
FILL FILL_37_DFFSR_39 ( );
FILL FILL_38_DFFSR_39 ( );
FILL FILL_39_DFFSR_39 ( );
FILL FILL_40_DFFSR_39 ( );
FILL FILL_41_DFFSR_39 ( );
FILL FILL_42_DFFSR_39 ( );
FILL FILL_43_DFFSR_39 ( );
FILL FILL_44_DFFSR_39 ( );
FILL FILL_45_DFFSR_39 ( );
FILL FILL_46_DFFSR_39 ( );
FILL FILL_47_DFFSR_39 ( );
FILL FILL_48_DFFSR_39 ( );
FILL FILL_49_DFFSR_39 ( );
FILL FILL_50_DFFSR_39 ( );
FILL FILL_51_DFFSR_39 ( );
FILL FILL_0_DFFSR_83 ( );
FILL FILL_1_DFFSR_83 ( );
FILL FILL_2_DFFSR_83 ( );
FILL FILL_3_DFFSR_83 ( );
FILL FILL_4_DFFSR_83 ( );
FILL FILL_5_DFFSR_83 ( );
FILL FILL_6_DFFSR_83 ( );
FILL FILL_7_DFFSR_83 ( );
FILL FILL_8_DFFSR_83 ( );
FILL FILL_9_DFFSR_83 ( );
FILL FILL_10_DFFSR_83 ( );
FILL FILL_11_DFFSR_83 ( );
FILL FILL_12_DFFSR_83 ( );
FILL FILL_13_DFFSR_83 ( );
FILL FILL_14_DFFSR_83 ( );
FILL FILL_15_DFFSR_83 ( );
FILL FILL_16_DFFSR_83 ( );
FILL FILL_17_DFFSR_83 ( );
FILL FILL_18_DFFSR_83 ( );
FILL FILL_19_DFFSR_83 ( );
FILL FILL_20_DFFSR_83 ( );
FILL FILL_21_DFFSR_83 ( );
FILL FILL_22_DFFSR_83 ( );
FILL FILL_23_DFFSR_83 ( );
FILL FILL_24_DFFSR_83 ( );
FILL FILL_25_DFFSR_83 ( );
FILL FILL_26_DFFSR_83 ( );
FILL FILL_27_DFFSR_83 ( );
FILL FILL_28_DFFSR_83 ( );
FILL FILL_29_DFFSR_83 ( );
FILL FILL_30_DFFSR_83 ( );
FILL FILL_31_DFFSR_83 ( );
FILL FILL_32_DFFSR_83 ( );
FILL FILL_33_DFFSR_83 ( );
FILL FILL_34_DFFSR_83 ( );
FILL FILL_35_DFFSR_83 ( );
FILL FILL_36_DFFSR_83 ( );
FILL FILL_37_DFFSR_83 ( );
FILL FILL_38_DFFSR_83 ( );
FILL FILL_39_DFFSR_83 ( );
FILL FILL_40_DFFSR_83 ( );
FILL FILL_41_DFFSR_83 ( );
FILL FILL_42_DFFSR_83 ( );
FILL FILL_43_DFFSR_83 ( );
FILL FILL_44_DFFSR_83 ( );
FILL FILL_45_DFFSR_83 ( );
FILL FILL_46_DFFSR_83 ( );
FILL FILL_47_DFFSR_83 ( );
FILL FILL_48_DFFSR_83 ( );
FILL FILL_49_DFFSR_83 ( );
FILL FILL_50_DFFSR_83 ( );
FILL FILL_51_DFFSR_83 ( );
FILL FILL_0_DFFSR_132 ( );
FILL FILL_1_DFFSR_132 ( );
FILL FILL_2_DFFSR_132 ( );
FILL FILL_3_DFFSR_132 ( );
FILL FILL_4_DFFSR_132 ( );
FILL FILL_5_DFFSR_132 ( );
FILL FILL_6_DFFSR_132 ( );
FILL FILL_7_DFFSR_132 ( );
FILL FILL_8_DFFSR_132 ( );
FILL FILL_9_DFFSR_132 ( );
FILL FILL_10_DFFSR_132 ( );
FILL FILL_11_DFFSR_132 ( );
FILL FILL_12_DFFSR_132 ( );
FILL FILL_13_DFFSR_132 ( );
FILL FILL_14_DFFSR_132 ( );
FILL FILL_15_DFFSR_132 ( );
FILL FILL_16_DFFSR_132 ( );
FILL FILL_17_DFFSR_132 ( );
FILL FILL_18_DFFSR_132 ( );
FILL FILL_19_DFFSR_132 ( );
FILL FILL_20_DFFSR_132 ( );
FILL FILL_21_DFFSR_132 ( );
FILL FILL_22_DFFSR_132 ( );
FILL FILL_23_DFFSR_132 ( );
FILL FILL_24_DFFSR_132 ( );
FILL FILL_25_DFFSR_132 ( );
FILL FILL_26_DFFSR_132 ( );
FILL FILL_27_DFFSR_132 ( );
FILL FILL_28_DFFSR_132 ( );
FILL FILL_29_DFFSR_132 ( );
FILL FILL_30_DFFSR_132 ( );
FILL FILL_31_DFFSR_132 ( );
FILL FILL_32_DFFSR_132 ( );
FILL FILL_33_DFFSR_132 ( );
FILL FILL_34_DFFSR_132 ( );
FILL FILL_35_DFFSR_132 ( );
FILL FILL_36_DFFSR_132 ( );
FILL FILL_37_DFFSR_132 ( );
FILL FILL_38_DFFSR_132 ( );
FILL FILL_39_DFFSR_132 ( );
FILL FILL_40_DFFSR_132 ( );
FILL FILL_41_DFFSR_132 ( );
FILL FILL_42_DFFSR_132 ( );
FILL FILL_43_DFFSR_132 ( );
FILL FILL_44_DFFSR_132 ( );
FILL FILL_45_DFFSR_132 ( );
FILL FILL_46_DFFSR_132 ( );
FILL FILL_47_DFFSR_132 ( );
FILL FILL_48_DFFSR_132 ( );
FILL FILL_49_DFFSR_132 ( );
FILL FILL_50_DFFSR_132 ( );
FILL FILL_0_NAND2X1_32 ( );
FILL FILL_1_NAND2X1_32 ( );
FILL FILL_2_NAND2X1_32 ( );
FILL FILL_3_NAND2X1_32 ( );
FILL FILL_4_NAND2X1_32 ( );
FILL FILL_5_NAND2X1_32 ( );
FILL FILL_6_NAND2X1_32 ( );
FILL FILL_0_NAND2X1_36 ( );
FILL FILL_1_NAND2X1_36 ( );
FILL FILL_2_NAND2X1_36 ( );
FILL FILL_3_NAND2X1_36 ( );
FILL FILL_4_NAND2X1_36 ( );
FILL FILL_5_NAND2X1_36 ( );
FILL FILL_6_NAND2X1_36 ( );
FILL FILL_0_DFFSR_205 ( );
FILL FILL_1_DFFSR_205 ( );
FILL FILL_2_DFFSR_205 ( );
FILL FILL_3_DFFSR_205 ( );
FILL FILL_4_DFFSR_205 ( );
FILL FILL_5_DFFSR_205 ( );
FILL FILL_6_DFFSR_205 ( );
FILL FILL_7_DFFSR_205 ( );
FILL FILL_8_DFFSR_205 ( );
FILL FILL_9_DFFSR_205 ( );
FILL FILL_10_DFFSR_205 ( );
FILL FILL_11_DFFSR_205 ( );
FILL FILL_12_DFFSR_205 ( );
FILL FILL_13_DFFSR_205 ( );
FILL FILL_14_DFFSR_205 ( );
FILL FILL_15_DFFSR_205 ( );
FILL FILL_16_DFFSR_205 ( );
FILL FILL_17_DFFSR_205 ( );
FILL FILL_18_DFFSR_205 ( );
FILL FILL_19_DFFSR_205 ( );
FILL FILL_20_DFFSR_205 ( );
FILL FILL_21_DFFSR_205 ( );
FILL FILL_22_DFFSR_205 ( );
FILL FILL_23_DFFSR_205 ( );
FILL FILL_24_DFFSR_205 ( );
FILL FILL_25_DFFSR_205 ( );
FILL FILL_26_DFFSR_205 ( );
FILL FILL_27_DFFSR_205 ( );
FILL FILL_28_DFFSR_205 ( );
FILL FILL_29_DFFSR_205 ( );
FILL FILL_30_DFFSR_205 ( );
FILL FILL_31_DFFSR_205 ( );
FILL FILL_32_DFFSR_205 ( );
FILL FILL_33_DFFSR_205 ( );
FILL FILL_34_DFFSR_205 ( );
FILL FILL_35_DFFSR_205 ( );
FILL FILL_36_DFFSR_205 ( );
FILL FILL_37_DFFSR_205 ( );
FILL FILL_38_DFFSR_205 ( );
FILL FILL_39_DFFSR_205 ( );
FILL FILL_40_DFFSR_205 ( );
FILL FILL_41_DFFSR_205 ( );
FILL FILL_42_DFFSR_205 ( );
FILL FILL_43_DFFSR_205 ( );
FILL FILL_44_DFFSR_205 ( );
FILL FILL_45_DFFSR_205 ( );
FILL FILL_46_DFFSR_205 ( );
FILL FILL_47_DFFSR_205 ( );
FILL FILL_48_DFFSR_205 ( );
FILL FILL_49_DFFSR_205 ( );
FILL FILL_50_DFFSR_205 ( );
FILL FILL_51_DFFSR_205 ( );
FILL FILL_0_OAI22X1_29 ( );
FILL FILL_1_OAI22X1_29 ( );
FILL FILL_2_OAI22X1_29 ( );
FILL FILL_3_OAI22X1_29 ( );
FILL FILL_4_OAI22X1_29 ( );
FILL FILL_5_OAI22X1_29 ( );
FILL FILL_6_OAI22X1_29 ( );
FILL FILL_7_OAI22X1_29 ( );
FILL FILL_8_OAI22X1_29 ( );
FILL FILL_9_OAI22X1_29 ( );
FILL FILL_10_OAI22X1_29 ( );
FILL FILL_0_NOR2X1_38 ( );
FILL FILL_1_NOR2X1_38 ( );
FILL FILL_2_NOR2X1_38 ( );
FILL FILL_3_NOR2X1_38 ( );
FILL FILL_4_NOR2X1_38 ( );
FILL FILL_5_NOR2X1_38 ( );
FILL FILL_6_NOR2X1_38 ( );
FILL FILL_0_NOR2X1_58 ( );
FILL FILL_1_NOR2X1_58 ( );
FILL FILL_2_NOR2X1_58 ( );
FILL FILL_3_NOR2X1_58 ( );
FILL FILL_4_NOR2X1_58 ( );
FILL FILL_5_NOR2X1_58 ( );
FILL FILL_6_NOR2X1_58 ( );
FILL FILL_0_OAI21X1_15 ( );
FILL FILL_1_OAI21X1_15 ( );
FILL FILL_2_OAI21X1_15 ( );
FILL FILL_3_OAI21X1_15 ( );
FILL FILL_4_OAI21X1_15 ( );
FILL FILL_5_OAI21X1_15 ( );
FILL FILL_6_OAI21X1_15 ( );
FILL FILL_7_OAI21X1_15 ( );
FILL FILL_8_OAI21X1_15 ( );
FILL FILL_9_OAI21X1_15 ( );
FILL FILL_0_NAND2X1_49 ( );
FILL FILL_1_NAND2X1_49 ( );
FILL FILL_2_NAND2X1_49 ( );
FILL FILL_3_NAND2X1_49 ( );
FILL FILL_4_NAND2X1_49 ( );
FILL FILL_5_NAND2X1_49 ( );
FILL FILL_6_NAND2X1_49 ( );
FILL FILL_0_DFFSR_181 ( );
FILL FILL_1_DFFSR_181 ( );
FILL FILL_2_DFFSR_181 ( );
FILL FILL_3_DFFSR_181 ( );
FILL FILL_4_DFFSR_181 ( );
FILL FILL_5_DFFSR_181 ( );
FILL FILL_6_DFFSR_181 ( );
FILL FILL_7_DFFSR_181 ( );
FILL FILL_8_DFFSR_181 ( );
FILL FILL_9_DFFSR_181 ( );
FILL FILL_10_DFFSR_181 ( );
FILL FILL_11_DFFSR_181 ( );
FILL FILL_12_DFFSR_181 ( );
FILL FILL_13_DFFSR_181 ( );
FILL FILL_14_DFFSR_181 ( );
FILL FILL_15_DFFSR_181 ( );
FILL FILL_16_DFFSR_181 ( );
FILL FILL_17_DFFSR_181 ( );
FILL FILL_18_DFFSR_181 ( );
FILL FILL_19_DFFSR_181 ( );
FILL FILL_20_DFFSR_181 ( );
FILL FILL_21_DFFSR_181 ( );
FILL FILL_22_DFFSR_181 ( );
FILL FILL_23_DFFSR_181 ( );
FILL FILL_24_DFFSR_181 ( );
FILL FILL_25_DFFSR_181 ( );
FILL FILL_26_DFFSR_181 ( );
FILL FILL_27_DFFSR_181 ( );
FILL FILL_28_DFFSR_181 ( );
FILL FILL_29_DFFSR_181 ( );
FILL FILL_30_DFFSR_181 ( );
FILL FILL_31_DFFSR_181 ( );
FILL FILL_32_DFFSR_181 ( );
FILL FILL_33_DFFSR_181 ( );
FILL FILL_34_DFFSR_181 ( );
FILL FILL_35_DFFSR_181 ( );
FILL FILL_36_DFFSR_181 ( );
FILL FILL_37_DFFSR_181 ( );
FILL FILL_38_DFFSR_181 ( );
FILL FILL_39_DFFSR_181 ( );
FILL FILL_40_DFFSR_181 ( );
FILL FILL_41_DFFSR_181 ( );
FILL FILL_42_DFFSR_181 ( );
FILL FILL_43_DFFSR_181 ( );
FILL FILL_44_DFFSR_181 ( );
FILL FILL_45_DFFSR_181 ( );
FILL FILL_46_DFFSR_181 ( );
FILL FILL_47_DFFSR_181 ( );
FILL FILL_48_DFFSR_181 ( );
FILL FILL_49_DFFSR_181 ( );
FILL FILL_50_DFFSR_181 ( );
FILL FILL_0_AND2X2_36 ( );
FILL FILL_1_AND2X2_36 ( );
FILL FILL_2_AND2X2_36 ( );
FILL FILL_3_AND2X2_36 ( );
FILL FILL_4_AND2X2_36 ( );
FILL FILL_5_AND2X2_36 ( );
FILL FILL_6_AND2X2_36 ( );
FILL FILL_7_AND2X2_36 ( );
FILL FILL_8_AND2X2_36 ( );
FILL FILL_0_NAND2X1_92 ( );
FILL FILL_1_NAND2X1_92 ( );
FILL FILL_2_NAND2X1_92 ( );
FILL FILL_3_NAND2X1_92 ( );
FILL FILL_4_NAND2X1_92 ( );
FILL FILL_5_NAND2X1_92 ( );
FILL FILL_6_NAND2X1_92 ( );
FILL FILL_0_NAND3X1_176 ( );
FILL FILL_1_NAND3X1_176 ( );
FILL FILL_2_NAND3X1_176 ( );
FILL FILL_3_NAND3X1_176 ( );
FILL FILL_4_NAND3X1_176 ( );
FILL FILL_5_NAND3X1_176 ( );
FILL FILL_6_NAND3X1_176 ( );
FILL FILL_7_NAND3X1_176 ( );
FILL FILL_8_NAND3X1_176 ( );
FILL FILL_9_NAND3X1_176 ( );
FILL FILL_0_NAND3X1_179 ( );
FILL FILL_1_NAND3X1_179 ( );
FILL FILL_2_NAND3X1_179 ( );
FILL FILL_3_NAND3X1_179 ( );
FILL FILL_4_NAND3X1_179 ( );
FILL FILL_5_NAND3X1_179 ( );
FILL FILL_6_NAND3X1_179 ( );
FILL FILL_7_NAND3X1_179 ( );
FILL FILL_8_NAND3X1_179 ( );
FILL FILL_0_AND2X2_33 ( );
FILL FILL_1_AND2X2_33 ( );
FILL FILL_2_AND2X2_33 ( );
FILL FILL_3_AND2X2_33 ( );
FILL FILL_4_AND2X2_33 ( );
FILL FILL_5_AND2X2_33 ( );
FILL FILL_6_AND2X2_33 ( );
FILL FILL_7_AND2X2_33 ( );
FILL FILL_8_AND2X2_33 ( );
FILL FILL_9_AND2X2_33 ( );
FILL FILL_0_NAND3X1_174 ( );
FILL FILL_1_NAND3X1_174 ( );
FILL FILL_2_NAND3X1_174 ( );
FILL FILL_3_NAND3X1_174 ( );
FILL FILL_4_NAND3X1_174 ( );
FILL FILL_5_NAND3X1_174 ( );
FILL FILL_6_NAND3X1_174 ( );
FILL FILL_7_NAND3X1_174 ( );
FILL FILL_8_NAND3X1_174 ( );
FILL FILL_0_AND2X2_31 ( );
FILL FILL_1_AND2X2_31 ( );
FILL FILL_2_AND2X2_31 ( );
FILL FILL_3_AND2X2_31 ( );
FILL FILL_4_AND2X2_31 ( );
FILL FILL_5_AND2X2_31 ( );
FILL FILL_6_AND2X2_31 ( );
FILL FILL_7_AND2X2_31 ( );
FILL FILL_8_AND2X2_31 ( );
FILL FILL_9_AND2X2_31 ( );
FILL FILL_0_AOI22X1_17 ( );
FILL FILL_1_AOI22X1_17 ( );
FILL FILL_2_AOI22X1_17 ( );
FILL FILL_3_AOI22X1_17 ( );
FILL FILL_4_AOI22X1_17 ( );
FILL FILL_5_AOI22X1_17 ( );
FILL FILL_6_AOI22X1_17 ( );
FILL FILL_7_AOI22X1_17 ( );
FILL FILL_8_AOI22X1_17 ( );
FILL FILL_9_AOI22X1_17 ( );
FILL FILL_10_AOI22X1_17 ( );
FILL FILL_0_AOI21X1_56 ( );
FILL FILL_1_AOI21X1_56 ( );
FILL FILL_2_AOI21X1_56 ( );
FILL FILL_3_AOI21X1_56 ( );
FILL FILL_4_AOI21X1_56 ( );
FILL FILL_5_AOI21X1_56 ( );
FILL FILL_6_AOI21X1_56 ( );
FILL FILL_7_AOI21X1_56 ( );
FILL FILL_8_AOI21X1_56 ( );
FILL FILL_9_AOI21X1_56 ( );
FILL FILL_0_NAND2X1_160 ( );
FILL FILL_1_NAND2X1_160 ( );
FILL FILL_2_NAND2X1_160 ( );
FILL FILL_3_NAND2X1_160 ( );
FILL FILL_4_NAND2X1_160 ( );
FILL FILL_5_NAND2X1_160 ( );
FILL FILL_6_NAND2X1_160 ( );
FILL FILL_0_NAND2X1_171 ( );
FILL FILL_1_NAND2X1_171 ( );
FILL FILL_2_NAND2X1_171 ( );
FILL FILL_3_NAND2X1_171 ( );
FILL FILL_4_NAND2X1_171 ( );
FILL FILL_5_NAND2X1_171 ( );
FILL FILL_6_NAND2X1_171 ( );
FILL FILL_0_NOR3X1_6 ( );
FILL FILL_1_NOR3X1_6 ( );
FILL FILL_2_NOR3X1_6 ( );
FILL FILL_3_NOR3X1_6 ( );
FILL FILL_4_NOR3X1_6 ( );
FILL FILL_5_NOR3X1_6 ( );
FILL FILL_6_NOR3X1_6 ( );
FILL FILL_7_NOR3X1_6 ( );
FILL FILL_8_NOR3X1_6 ( );
FILL FILL_9_NOR3X1_6 ( );
FILL FILL_10_NOR3X1_6 ( );
FILL FILL_11_NOR3X1_6 ( );
FILL FILL_12_NOR3X1_6 ( );
FILL FILL_13_NOR3X1_6 ( );
FILL FILL_14_NOR3X1_6 ( );
FILL FILL_15_NOR3X1_6 ( );
FILL FILL_16_NOR3X1_6 ( );
FILL FILL_17_NOR3X1_6 ( );
FILL FILL_18_NOR3X1_6 ( );
FILL FILL_0_OAI21X1_109 ( );
FILL FILL_1_OAI21X1_109 ( );
FILL FILL_2_OAI21X1_109 ( );
FILL FILL_3_OAI21X1_109 ( );
FILL FILL_4_OAI21X1_109 ( );
FILL FILL_5_OAI21X1_109 ( );
FILL FILL_6_OAI21X1_109 ( );
FILL FILL_7_OAI21X1_109 ( );
FILL FILL_8_OAI21X1_109 ( );
FILL FILL_0_NAND3X1_247 ( );
FILL FILL_1_NAND3X1_247 ( );
FILL FILL_2_NAND3X1_247 ( );
FILL FILL_3_NAND3X1_247 ( );
FILL FILL_4_NAND3X1_247 ( );
FILL FILL_5_NAND3X1_247 ( );
FILL FILL_6_NAND3X1_247 ( );
FILL FILL_7_NAND3X1_247 ( );
FILL FILL_8_NAND3X1_247 ( );
FILL FILL_0_INVX1_210 ( );
FILL FILL_1_INVX1_210 ( );
FILL FILL_2_INVX1_210 ( );
FILL FILL_3_INVX1_210 ( );
FILL FILL_4_INVX1_210 ( );
FILL FILL_0_DFFSR_79 ( );
FILL FILL_1_DFFSR_79 ( );
FILL FILL_2_DFFSR_79 ( );
FILL FILL_3_DFFSR_79 ( );
FILL FILL_4_DFFSR_79 ( );
FILL FILL_5_DFFSR_79 ( );
FILL FILL_6_DFFSR_79 ( );
FILL FILL_7_DFFSR_79 ( );
FILL FILL_8_DFFSR_79 ( );
FILL FILL_9_DFFSR_79 ( );
FILL FILL_10_DFFSR_79 ( );
FILL FILL_11_DFFSR_79 ( );
FILL FILL_12_DFFSR_79 ( );
FILL FILL_13_DFFSR_79 ( );
FILL FILL_14_DFFSR_79 ( );
FILL FILL_15_DFFSR_79 ( );
FILL FILL_16_DFFSR_79 ( );
FILL FILL_17_DFFSR_79 ( );
FILL FILL_18_DFFSR_79 ( );
FILL FILL_19_DFFSR_79 ( );
FILL FILL_20_DFFSR_79 ( );
FILL FILL_21_DFFSR_79 ( );
FILL FILL_22_DFFSR_79 ( );
FILL FILL_23_DFFSR_79 ( );
FILL FILL_24_DFFSR_79 ( );
FILL FILL_25_DFFSR_79 ( );
FILL FILL_26_DFFSR_79 ( );
FILL FILL_27_DFFSR_79 ( );
FILL FILL_28_DFFSR_79 ( );
FILL FILL_29_DFFSR_79 ( );
FILL FILL_30_DFFSR_79 ( );
FILL FILL_31_DFFSR_79 ( );
FILL FILL_32_DFFSR_79 ( );
FILL FILL_33_DFFSR_79 ( );
FILL FILL_34_DFFSR_79 ( );
FILL FILL_35_DFFSR_79 ( );
FILL FILL_36_DFFSR_79 ( );
FILL FILL_37_DFFSR_79 ( );
FILL FILL_38_DFFSR_79 ( );
FILL FILL_39_DFFSR_79 ( );
FILL FILL_40_DFFSR_79 ( );
FILL FILL_41_DFFSR_79 ( );
FILL FILL_42_DFFSR_79 ( );
FILL FILL_43_DFFSR_79 ( );
FILL FILL_44_DFFSR_79 ( );
FILL FILL_45_DFFSR_79 ( );
FILL FILL_46_DFFSR_79 ( );
FILL FILL_47_DFFSR_79 ( );
FILL FILL_48_DFFSR_79 ( );
FILL FILL_49_DFFSR_79 ( );
FILL FILL_50_DFFSR_79 ( );
FILL FILL_0_XOR2X1_9 ( );
FILL FILL_1_XOR2X1_9 ( );
FILL FILL_2_XOR2X1_9 ( );
FILL FILL_3_XOR2X1_9 ( );
FILL FILL_4_XOR2X1_9 ( );
FILL FILL_5_XOR2X1_9 ( );
FILL FILL_6_XOR2X1_9 ( );
FILL FILL_7_XOR2X1_9 ( );
FILL FILL_8_XOR2X1_9 ( );
FILL FILL_9_XOR2X1_9 ( );
FILL FILL_10_XOR2X1_9 ( );
FILL FILL_11_XOR2X1_9 ( );
FILL FILL_12_XOR2X1_9 ( );
FILL FILL_13_XOR2X1_9 ( );
FILL FILL_14_XOR2X1_9 ( );
FILL FILL_15_XOR2X1_9 ( );
FILL FILL_0_NAND2X1_173 ( );
FILL FILL_1_NAND2X1_173 ( );
FILL FILL_2_NAND2X1_173 ( );
FILL FILL_3_NAND2X1_173 ( );
FILL FILL_4_NAND2X1_173 ( );
FILL FILL_5_NAND2X1_173 ( );
FILL FILL_6_NAND2X1_173 ( );
FILL FILL_0_OAI21X1_113 ( );
FILL FILL_1_OAI21X1_113 ( );
FILL FILL_2_OAI21X1_113 ( );
FILL FILL_3_OAI21X1_113 ( );
FILL FILL_4_OAI21X1_113 ( );
FILL FILL_5_OAI21X1_113 ( );
FILL FILL_6_OAI21X1_113 ( );
FILL FILL_7_OAI21X1_113 ( );
FILL FILL_8_OAI21X1_113 ( );
FILL FILL_0_INVX1_20 ( );
FILL FILL_1_INVX1_20 ( );
FILL FILL_2_INVX1_20 ( );
FILL FILL_3_INVX1_20 ( );
FILL FILL_0_CLKBUF1_8 ( );
FILL FILL_1_CLKBUF1_8 ( );
FILL FILL_2_CLKBUF1_8 ( );
FILL FILL_3_CLKBUF1_8 ( );
FILL FILL_4_CLKBUF1_8 ( );
FILL FILL_5_CLKBUF1_8 ( );
FILL FILL_6_CLKBUF1_8 ( );
FILL FILL_7_CLKBUF1_8 ( );
FILL FILL_8_CLKBUF1_8 ( );
FILL FILL_9_CLKBUF1_8 ( );
FILL FILL_10_CLKBUF1_8 ( );
FILL FILL_11_CLKBUF1_8 ( );
FILL FILL_12_CLKBUF1_8 ( );
FILL FILL_13_CLKBUF1_8 ( );
FILL FILL_14_CLKBUF1_8 ( );
FILL FILL_15_CLKBUF1_8 ( );
FILL FILL_16_CLKBUF1_8 ( );
FILL FILL_17_CLKBUF1_8 ( );
FILL FILL_18_CLKBUF1_8 ( );
FILL FILL_19_CLKBUF1_8 ( );
FILL FILL_20_CLKBUF1_8 ( );
FILL FILL_0_INVX1_58 ( );
FILL FILL_1_INVX1_58 ( );
FILL FILL_2_INVX1_58 ( );
FILL FILL_3_INVX1_58 ( );
FILL FILL_4_INVX1_58 ( );
FILL FILL_0_CLKBUF1_36 ( );
FILL FILL_1_CLKBUF1_36 ( );
FILL FILL_2_CLKBUF1_36 ( );
FILL FILL_3_CLKBUF1_36 ( );
FILL FILL_4_CLKBUF1_36 ( );
FILL FILL_5_CLKBUF1_36 ( );
FILL FILL_6_CLKBUF1_36 ( );
FILL FILL_7_CLKBUF1_36 ( );
FILL FILL_8_CLKBUF1_36 ( );
FILL FILL_9_CLKBUF1_36 ( );
FILL FILL_10_CLKBUF1_36 ( );
FILL FILL_11_CLKBUF1_36 ( );
FILL FILL_12_CLKBUF1_36 ( );
FILL FILL_13_CLKBUF1_36 ( );
FILL FILL_14_CLKBUF1_36 ( );
FILL FILL_15_CLKBUF1_36 ( );
FILL FILL_16_CLKBUF1_36 ( );
FILL FILL_17_CLKBUF1_36 ( );
FILL FILL_18_CLKBUF1_36 ( );
FILL FILL_19_CLKBUF1_36 ( );
FILL FILL_20_CLKBUF1_36 ( );
FILL FILL_0_OAI22X1_2 ( );
FILL FILL_1_OAI22X1_2 ( );
FILL FILL_2_OAI22X1_2 ( );
FILL FILL_3_OAI22X1_2 ( );
FILL FILL_4_OAI22X1_2 ( );
FILL FILL_5_OAI22X1_2 ( );
FILL FILL_6_OAI22X1_2 ( );
FILL FILL_7_OAI22X1_2 ( );
FILL FILL_8_OAI22X1_2 ( );
FILL FILL_9_OAI22X1_2 ( );
FILL FILL_10_OAI22X1_2 ( );
FILL FILL_0_DFFSR_131 ( );
FILL FILL_1_DFFSR_131 ( );
FILL FILL_2_DFFSR_131 ( );
FILL FILL_3_DFFSR_131 ( );
FILL FILL_4_DFFSR_131 ( );
FILL FILL_5_DFFSR_131 ( );
FILL FILL_6_DFFSR_131 ( );
FILL FILL_7_DFFSR_131 ( );
FILL FILL_8_DFFSR_131 ( );
FILL FILL_9_DFFSR_131 ( );
FILL FILL_10_DFFSR_131 ( );
FILL FILL_11_DFFSR_131 ( );
FILL FILL_12_DFFSR_131 ( );
FILL FILL_13_DFFSR_131 ( );
FILL FILL_14_DFFSR_131 ( );
FILL FILL_15_DFFSR_131 ( );
FILL FILL_16_DFFSR_131 ( );
FILL FILL_17_DFFSR_131 ( );
FILL FILL_18_DFFSR_131 ( );
FILL FILL_19_DFFSR_131 ( );
FILL FILL_20_DFFSR_131 ( );
FILL FILL_21_DFFSR_131 ( );
FILL FILL_22_DFFSR_131 ( );
FILL FILL_23_DFFSR_131 ( );
FILL FILL_24_DFFSR_131 ( );
FILL FILL_25_DFFSR_131 ( );
FILL FILL_26_DFFSR_131 ( );
FILL FILL_27_DFFSR_131 ( );
FILL FILL_28_DFFSR_131 ( );
FILL FILL_29_DFFSR_131 ( );
FILL FILL_30_DFFSR_131 ( );
FILL FILL_31_DFFSR_131 ( );
FILL FILL_32_DFFSR_131 ( );
FILL FILL_33_DFFSR_131 ( );
FILL FILL_34_DFFSR_131 ( );
FILL FILL_35_DFFSR_131 ( );
FILL FILL_36_DFFSR_131 ( );
FILL FILL_37_DFFSR_131 ( );
FILL FILL_38_DFFSR_131 ( );
FILL FILL_39_DFFSR_131 ( );
FILL FILL_40_DFFSR_131 ( );
FILL FILL_41_DFFSR_131 ( );
FILL FILL_42_DFFSR_131 ( );
FILL FILL_43_DFFSR_131 ( );
FILL FILL_44_DFFSR_131 ( );
FILL FILL_45_DFFSR_131 ( );
FILL FILL_46_DFFSR_131 ( );
FILL FILL_47_DFFSR_131 ( );
FILL FILL_48_DFFSR_131 ( );
FILL FILL_49_DFFSR_131 ( );
FILL FILL_50_DFFSR_131 ( );
FILL FILL_51_DFFSR_131 ( );
FILL FILL_0_DFFSR_136 ( );
FILL FILL_1_DFFSR_136 ( );
FILL FILL_2_DFFSR_136 ( );
FILL FILL_3_DFFSR_136 ( );
FILL FILL_4_DFFSR_136 ( );
FILL FILL_5_DFFSR_136 ( );
FILL FILL_6_DFFSR_136 ( );
FILL FILL_7_DFFSR_136 ( );
FILL FILL_8_DFFSR_136 ( );
FILL FILL_9_DFFSR_136 ( );
FILL FILL_10_DFFSR_136 ( );
FILL FILL_11_DFFSR_136 ( );
FILL FILL_12_DFFSR_136 ( );
FILL FILL_13_DFFSR_136 ( );
FILL FILL_14_DFFSR_136 ( );
FILL FILL_15_DFFSR_136 ( );
FILL FILL_16_DFFSR_136 ( );
FILL FILL_17_DFFSR_136 ( );
FILL FILL_18_DFFSR_136 ( );
FILL FILL_19_DFFSR_136 ( );
FILL FILL_20_DFFSR_136 ( );
FILL FILL_21_DFFSR_136 ( );
FILL FILL_22_DFFSR_136 ( );
FILL FILL_23_DFFSR_136 ( );
FILL FILL_24_DFFSR_136 ( );
FILL FILL_25_DFFSR_136 ( );
FILL FILL_26_DFFSR_136 ( );
FILL FILL_27_DFFSR_136 ( );
FILL FILL_28_DFFSR_136 ( );
FILL FILL_29_DFFSR_136 ( );
FILL FILL_30_DFFSR_136 ( );
FILL FILL_31_DFFSR_136 ( );
FILL FILL_32_DFFSR_136 ( );
FILL FILL_33_DFFSR_136 ( );
FILL FILL_34_DFFSR_136 ( );
FILL FILL_35_DFFSR_136 ( );
FILL FILL_36_DFFSR_136 ( );
FILL FILL_37_DFFSR_136 ( );
FILL FILL_38_DFFSR_136 ( );
FILL FILL_39_DFFSR_136 ( );
FILL FILL_40_DFFSR_136 ( );
FILL FILL_41_DFFSR_136 ( );
FILL FILL_42_DFFSR_136 ( );
FILL FILL_43_DFFSR_136 ( );
FILL FILL_44_DFFSR_136 ( );
FILL FILL_45_DFFSR_136 ( );
FILL FILL_46_DFFSR_136 ( );
FILL FILL_47_DFFSR_136 ( );
FILL FILL_48_DFFSR_136 ( );
FILL FILL_49_DFFSR_136 ( );
FILL FILL_50_DFFSR_136 ( );
FILL FILL_0_INVX1_72 ( );
FILL FILL_1_INVX1_72 ( );
FILL FILL_2_INVX1_72 ( );
FILL FILL_3_INVX1_72 ( );
FILL FILL_4_INVX1_72 ( );
FILL FILL_0_NAND3X1_128 ( );
FILL FILL_1_NAND3X1_128 ( );
FILL FILL_2_NAND3X1_128 ( );
FILL FILL_3_NAND3X1_128 ( );
FILL FILL_4_NAND3X1_128 ( );
FILL FILL_5_NAND3X1_128 ( );
FILL FILL_6_NAND3X1_128 ( );
FILL FILL_7_NAND3X1_128 ( );
FILL FILL_8_NAND3X1_128 ( );
FILL FILL_0_NAND3X1_78 ( );
FILL FILL_1_NAND3X1_78 ( );
FILL FILL_2_NAND3X1_78 ( );
FILL FILL_3_NAND3X1_78 ( );
FILL FILL_4_NAND3X1_78 ( );
FILL FILL_5_NAND3X1_78 ( );
FILL FILL_6_NAND3X1_78 ( );
FILL FILL_7_NAND3X1_78 ( );
FILL FILL_8_NAND3X1_78 ( );
FILL FILL_9_NAND3X1_78 ( );
FILL FILL_0_INVX1_70 ( );
FILL FILL_1_INVX1_70 ( );
FILL FILL_2_INVX1_70 ( );
FILL FILL_3_INVX1_70 ( );
FILL FILL_4_INVX1_70 ( );
FILL FILL_0_INVX1_90 ( );
FILL FILL_1_INVX1_90 ( );
FILL FILL_2_INVX1_90 ( );
FILL FILL_3_INVX1_90 ( );
FILL FILL_4_INVX1_90 ( );
FILL FILL_0_DFFSR_178 ( );
FILL FILL_1_DFFSR_178 ( );
FILL FILL_2_DFFSR_178 ( );
FILL FILL_3_DFFSR_178 ( );
FILL FILL_4_DFFSR_178 ( );
FILL FILL_5_DFFSR_178 ( );
FILL FILL_6_DFFSR_178 ( );
FILL FILL_7_DFFSR_178 ( );
FILL FILL_8_DFFSR_178 ( );
FILL FILL_9_DFFSR_178 ( );
FILL FILL_10_DFFSR_178 ( );
FILL FILL_11_DFFSR_178 ( );
FILL FILL_12_DFFSR_178 ( );
FILL FILL_13_DFFSR_178 ( );
FILL FILL_14_DFFSR_178 ( );
FILL FILL_15_DFFSR_178 ( );
FILL FILL_16_DFFSR_178 ( );
FILL FILL_17_DFFSR_178 ( );
FILL FILL_18_DFFSR_178 ( );
FILL FILL_19_DFFSR_178 ( );
FILL FILL_20_DFFSR_178 ( );
FILL FILL_21_DFFSR_178 ( );
FILL FILL_22_DFFSR_178 ( );
FILL FILL_23_DFFSR_178 ( );
FILL FILL_24_DFFSR_178 ( );
FILL FILL_25_DFFSR_178 ( );
FILL FILL_26_DFFSR_178 ( );
FILL FILL_27_DFFSR_178 ( );
FILL FILL_28_DFFSR_178 ( );
FILL FILL_29_DFFSR_178 ( );
FILL FILL_30_DFFSR_178 ( );
FILL FILL_31_DFFSR_178 ( );
FILL FILL_32_DFFSR_178 ( );
FILL FILL_33_DFFSR_178 ( );
FILL FILL_34_DFFSR_178 ( );
FILL FILL_35_DFFSR_178 ( );
FILL FILL_36_DFFSR_178 ( );
FILL FILL_37_DFFSR_178 ( );
FILL FILL_38_DFFSR_178 ( );
FILL FILL_39_DFFSR_178 ( );
FILL FILL_40_DFFSR_178 ( );
FILL FILL_41_DFFSR_178 ( );
FILL FILL_42_DFFSR_178 ( );
FILL FILL_43_DFFSR_178 ( );
FILL FILL_44_DFFSR_178 ( );
FILL FILL_45_DFFSR_178 ( );
FILL FILL_46_DFFSR_178 ( );
FILL FILL_47_DFFSR_178 ( );
FILL FILL_48_DFFSR_178 ( );
FILL FILL_49_DFFSR_178 ( );
FILL FILL_50_DFFSR_178 ( );
FILL FILL_0_NAND2X1_118 ( );
FILL FILL_1_NAND2X1_118 ( );
FILL FILL_2_NAND2X1_118 ( );
FILL FILL_3_NAND2X1_118 ( );
FILL FILL_4_NAND2X1_118 ( );
FILL FILL_5_NAND2X1_118 ( );
FILL FILL_6_NAND2X1_118 ( );
FILL FILL_0_INVX1_166 ( );
FILL FILL_1_INVX1_166 ( );
FILL FILL_2_INVX1_166 ( );
FILL FILL_3_INVX1_166 ( );
FILL FILL_4_INVX1_166 ( );
FILL FILL_0_NAND2X1_110 ( );
FILL FILL_1_NAND2X1_110 ( );
FILL FILL_2_NAND2X1_110 ( );
FILL FILL_3_NAND2X1_110 ( );
FILL FILL_4_NAND2X1_110 ( );
FILL FILL_5_NAND2X1_110 ( );
FILL FILL_6_NAND2X1_110 ( );
FILL FILL_0_NAND2X1_84 ( );
FILL FILL_1_NAND2X1_84 ( );
FILL FILL_2_NAND2X1_84 ( );
FILL FILL_3_NAND2X1_84 ( );
FILL FILL_4_NAND2X1_84 ( );
FILL FILL_5_NAND2X1_84 ( );
FILL FILL_6_NAND2X1_84 ( );
FILL FILL_0_NAND3X1_178 ( );
FILL FILL_1_NAND3X1_178 ( );
FILL FILL_2_NAND3X1_178 ( );
FILL FILL_3_NAND3X1_178 ( );
FILL FILL_4_NAND3X1_178 ( );
FILL FILL_5_NAND3X1_178 ( );
FILL FILL_6_NAND3X1_178 ( );
FILL FILL_7_NAND3X1_178 ( );
FILL FILL_8_NAND3X1_178 ( );
FILL FILL_9_NAND3X1_178 ( );
FILL FILL_0_NAND3X1_175 ( );
FILL FILL_1_NAND3X1_175 ( );
FILL FILL_2_NAND3X1_175 ( );
FILL FILL_3_NAND3X1_175 ( );
FILL FILL_4_NAND3X1_175 ( );
FILL FILL_5_NAND3X1_175 ( );
FILL FILL_6_NAND3X1_175 ( );
FILL FILL_7_NAND3X1_175 ( );
FILL FILL_8_NAND3X1_175 ( );
FILL FILL_0_NAND2X1_85 ( );
FILL FILL_1_NAND2X1_85 ( );
FILL FILL_2_NAND2X1_85 ( );
FILL FILL_3_NAND2X1_85 ( );
FILL FILL_4_NAND2X1_85 ( );
FILL FILL_5_NAND2X1_85 ( );
FILL FILL_6_NAND2X1_85 ( );
FILL FILL_0_NAND2X1_86 ( );
FILL FILL_1_NAND2X1_86 ( );
FILL FILL_2_NAND2X1_86 ( );
FILL FILL_3_NAND2X1_86 ( );
FILL FILL_4_NAND2X1_86 ( );
FILL FILL_5_NAND2X1_86 ( );
FILL FILL_6_NAND2X1_86 ( );
FILL FILL_0_NAND2X1_87 ( );
FILL FILL_1_NAND2X1_87 ( );
FILL FILL_2_NAND2X1_87 ( );
FILL FILL_3_NAND2X1_87 ( );
FILL FILL_4_NAND2X1_87 ( );
FILL FILL_5_NAND2X1_87 ( );
FILL FILL_6_NAND2X1_87 ( );
FILL FILL_0_INVX1_132 ( );
FILL FILL_1_INVX1_132 ( );
FILL FILL_2_INVX1_132 ( );
FILL FILL_3_INVX1_132 ( );
FILL FILL_0_DFFPOSX1_23 ( );
FILL FILL_1_DFFPOSX1_23 ( );
FILL FILL_2_DFFPOSX1_23 ( );
FILL FILL_3_DFFPOSX1_23 ( );
FILL FILL_4_DFFPOSX1_23 ( );
FILL FILL_5_DFFPOSX1_23 ( );
FILL FILL_6_DFFPOSX1_23 ( );
FILL FILL_7_DFFPOSX1_23 ( );
FILL FILL_8_DFFPOSX1_23 ( );
FILL FILL_9_DFFPOSX1_23 ( );
FILL FILL_10_DFFPOSX1_23 ( );
FILL FILL_11_DFFPOSX1_23 ( );
FILL FILL_12_DFFPOSX1_23 ( );
FILL FILL_13_DFFPOSX1_23 ( );
FILL FILL_14_DFFPOSX1_23 ( );
FILL FILL_15_DFFPOSX1_23 ( );
FILL FILL_16_DFFPOSX1_23 ( );
FILL FILL_17_DFFPOSX1_23 ( );
FILL FILL_18_DFFPOSX1_23 ( );
FILL FILL_19_DFFPOSX1_23 ( );
FILL FILL_20_DFFPOSX1_23 ( );
FILL FILL_21_DFFPOSX1_23 ( );
FILL FILL_22_DFFPOSX1_23 ( );
FILL FILL_23_DFFPOSX1_23 ( );
FILL FILL_24_DFFPOSX1_23 ( );
FILL FILL_25_DFFPOSX1_23 ( );
FILL FILL_26_DFFPOSX1_23 ( );
FILL FILL_27_DFFPOSX1_23 ( );
FILL FILL_0_INVX1_209 ( );
FILL FILL_1_INVX1_209 ( );
FILL FILL_2_INVX1_209 ( );
FILL FILL_3_INVX1_209 ( );
FILL FILL_4_INVX1_209 ( );
FILL FILL_0_AOI21X1_63 ( );
FILL FILL_1_AOI21X1_63 ( );
FILL FILL_2_AOI21X1_63 ( );
FILL FILL_3_AOI21X1_63 ( );
FILL FILL_4_AOI21X1_63 ( );
FILL FILL_5_AOI21X1_63 ( );
FILL FILL_6_AOI21X1_63 ( );
FILL FILL_7_AOI21X1_63 ( );
FILL FILL_8_AOI21X1_63 ( );
FILL FILL_0_NAND2X1_157 ( );
FILL FILL_1_NAND2X1_157 ( );
FILL FILL_2_NAND2X1_157 ( );
FILL FILL_3_NAND2X1_157 ( );
FILL FILL_4_NAND2X1_157 ( );
FILL FILL_5_NAND2X1_157 ( );
FILL FILL_6_NAND2X1_157 ( );
FILL FILL_0_OAI21X1_110 ( );
FILL FILL_1_OAI21X1_110 ( );
FILL FILL_2_OAI21X1_110 ( );
FILL FILL_3_OAI21X1_110 ( );
FILL FILL_4_OAI21X1_110 ( );
FILL FILL_5_OAI21X1_110 ( );
FILL FILL_6_OAI21X1_110 ( );
FILL FILL_7_OAI21X1_110 ( );
FILL FILL_8_OAI21X1_110 ( );
FILL FILL_0_DFFSR_18 ( );
FILL FILL_1_DFFSR_18 ( );
FILL FILL_2_DFFSR_18 ( );
FILL FILL_3_DFFSR_18 ( );
FILL FILL_4_DFFSR_18 ( );
FILL FILL_5_DFFSR_18 ( );
FILL FILL_6_DFFSR_18 ( );
FILL FILL_7_DFFSR_18 ( );
FILL FILL_8_DFFSR_18 ( );
FILL FILL_9_DFFSR_18 ( );
FILL FILL_10_DFFSR_18 ( );
FILL FILL_11_DFFSR_18 ( );
FILL FILL_12_DFFSR_18 ( );
FILL FILL_13_DFFSR_18 ( );
FILL FILL_14_DFFSR_18 ( );
FILL FILL_15_DFFSR_18 ( );
FILL FILL_16_DFFSR_18 ( );
FILL FILL_17_DFFSR_18 ( );
FILL FILL_18_DFFSR_18 ( );
FILL FILL_19_DFFSR_18 ( );
FILL FILL_20_DFFSR_18 ( );
FILL FILL_21_DFFSR_18 ( );
FILL FILL_22_DFFSR_18 ( );
FILL FILL_23_DFFSR_18 ( );
FILL FILL_24_DFFSR_18 ( );
FILL FILL_25_DFFSR_18 ( );
FILL FILL_26_DFFSR_18 ( );
FILL FILL_27_DFFSR_18 ( );
FILL FILL_28_DFFSR_18 ( );
FILL FILL_29_DFFSR_18 ( );
FILL FILL_30_DFFSR_18 ( );
FILL FILL_31_DFFSR_18 ( );
FILL FILL_32_DFFSR_18 ( );
FILL FILL_33_DFFSR_18 ( );
FILL FILL_34_DFFSR_18 ( );
FILL FILL_35_DFFSR_18 ( );
FILL FILL_36_DFFSR_18 ( );
FILL FILL_37_DFFSR_18 ( );
FILL FILL_38_DFFSR_18 ( );
FILL FILL_39_DFFSR_18 ( );
FILL FILL_40_DFFSR_18 ( );
FILL FILL_41_DFFSR_18 ( );
FILL FILL_42_DFFSR_18 ( );
FILL FILL_43_DFFSR_18 ( );
FILL FILL_44_DFFSR_18 ( );
FILL FILL_45_DFFSR_18 ( );
FILL FILL_46_DFFSR_18 ( );
FILL FILL_47_DFFSR_18 ( );
FILL FILL_48_DFFSR_18 ( );
FILL FILL_49_DFFSR_18 ( );
FILL FILL_50_DFFSR_18 ( );
FILL FILL_0_NOR2X1_80 ( );
FILL FILL_1_NOR2X1_80 ( );
FILL FILL_2_NOR2X1_80 ( );
FILL FILL_3_NOR2X1_80 ( );
FILL FILL_4_NOR2X1_80 ( );
FILL FILL_5_NOR2X1_80 ( );
FILL FILL_6_NOR2X1_80 ( );
FILL FILL_0_AOI21X1_66 ( );
FILL FILL_1_AOI21X1_66 ( );
FILL FILL_2_AOI21X1_66 ( );
FILL FILL_3_AOI21X1_66 ( );
FILL FILL_4_AOI21X1_66 ( );
FILL FILL_5_AOI21X1_66 ( );
FILL FILL_6_AOI21X1_66 ( );
FILL FILL_7_AOI21X1_66 ( );
FILL FILL_8_AOI21X1_66 ( );
FILL FILL_0_AOI21X1_67 ( );
FILL FILL_1_AOI21X1_67 ( );
FILL FILL_2_AOI21X1_67 ( );
FILL FILL_3_AOI21X1_67 ( );
FILL FILL_4_AOI21X1_67 ( );
FILL FILL_5_AOI21X1_67 ( );
FILL FILL_6_AOI21X1_67 ( );
FILL FILL_7_AOI21X1_67 ( );
FILL FILL_8_AOI21X1_67 ( );
FILL FILL_0_OAI21X1_115 ( );
FILL FILL_1_OAI21X1_115 ( );
FILL FILL_2_OAI21X1_115 ( );
FILL FILL_3_OAI21X1_115 ( );
FILL FILL_4_OAI21X1_115 ( );
FILL FILL_5_OAI21X1_115 ( );
FILL FILL_6_OAI21X1_115 ( );
FILL FILL_7_OAI21X1_115 ( );
FILL FILL_8_OAI21X1_115 ( );
FILL FILL_0_INVX1_215 ( );
FILL FILL_1_INVX1_215 ( );
FILL FILL_2_INVX1_215 ( );
FILL FILL_3_INVX1_215 ( );
FILL FILL_4_INVX1_215 ( );
FILL FILL_0_NOR2X1_78 ( );
FILL FILL_1_NOR2X1_78 ( );
FILL FILL_2_NOR2X1_78 ( );
FILL FILL_3_NOR2X1_78 ( );
FILL FILL_4_NOR2X1_78 ( );
FILL FILL_5_NOR2X1_78 ( );
FILL FILL_6_NOR2X1_78 ( );
FILL FILL_0_OAI22X1_8 ( );
FILL FILL_1_OAI22X1_8 ( );
FILL FILL_2_OAI22X1_8 ( );
FILL FILL_3_OAI22X1_8 ( );
FILL FILL_4_OAI22X1_8 ( );
FILL FILL_5_OAI22X1_8 ( );
FILL FILL_6_OAI22X1_8 ( );
FILL FILL_7_OAI22X1_8 ( );
FILL FILL_8_OAI22X1_8 ( );
FILL FILL_9_OAI22X1_8 ( );
FILL FILL_10_OAI22X1_8 ( );
FILL FILL_11_OAI22X1_8 ( );
FILL FILL_0_INVX1_19 ( );
FILL FILL_1_INVX1_19 ( );
FILL FILL_2_INVX1_19 ( );
FILL FILL_3_INVX1_19 ( );
FILL FILL_4_INVX1_19 ( );
FILL FILL_0_DFFSR_128 ( );
FILL FILL_1_DFFSR_128 ( );
FILL FILL_2_DFFSR_128 ( );
FILL FILL_3_DFFSR_128 ( );
FILL FILL_4_DFFSR_128 ( );
FILL FILL_5_DFFSR_128 ( );
FILL FILL_6_DFFSR_128 ( );
FILL FILL_7_DFFSR_128 ( );
FILL FILL_8_DFFSR_128 ( );
FILL FILL_9_DFFSR_128 ( );
FILL FILL_10_DFFSR_128 ( );
FILL FILL_11_DFFSR_128 ( );
FILL FILL_12_DFFSR_128 ( );
FILL FILL_13_DFFSR_128 ( );
FILL FILL_14_DFFSR_128 ( );
FILL FILL_15_DFFSR_128 ( );
FILL FILL_16_DFFSR_128 ( );
FILL FILL_17_DFFSR_128 ( );
FILL FILL_18_DFFSR_128 ( );
FILL FILL_19_DFFSR_128 ( );
FILL FILL_20_DFFSR_128 ( );
FILL FILL_21_DFFSR_128 ( );
FILL FILL_22_DFFSR_128 ( );
FILL FILL_23_DFFSR_128 ( );
FILL FILL_24_DFFSR_128 ( );
FILL FILL_25_DFFSR_128 ( );
FILL FILL_26_DFFSR_128 ( );
FILL FILL_27_DFFSR_128 ( );
FILL FILL_28_DFFSR_128 ( );
FILL FILL_29_DFFSR_128 ( );
FILL FILL_30_DFFSR_128 ( );
FILL FILL_31_DFFSR_128 ( );
FILL FILL_32_DFFSR_128 ( );
FILL FILL_33_DFFSR_128 ( );
FILL FILL_34_DFFSR_128 ( );
FILL FILL_35_DFFSR_128 ( );
FILL FILL_36_DFFSR_128 ( );
FILL FILL_37_DFFSR_128 ( );
FILL FILL_38_DFFSR_128 ( );
FILL FILL_39_DFFSR_128 ( );
FILL FILL_40_DFFSR_128 ( );
FILL FILL_41_DFFSR_128 ( );
FILL FILL_42_DFFSR_128 ( );
FILL FILL_43_DFFSR_128 ( );
FILL FILL_44_DFFSR_128 ( );
FILL FILL_45_DFFSR_128 ( );
FILL FILL_46_DFFSR_128 ( );
FILL FILL_47_DFFSR_128 ( );
FILL FILL_48_DFFSR_128 ( );
FILL FILL_49_DFFSR_128 ( );
FILL FILL_50_DFFSR_128 ( );
FILL FILL_0_AND2X2_16 ( );
FILL FILL_1_AND2X2_16 ( );
FILL FILL_2_AND2X2_16 ( );
FILL FILL_3_AND2X2_16 ( );
FILL FILL_4_AND2X2_16 ( );
FILL FILL_5_AND2X2_16 ( );
FILL FILL_6_AND2X2_16 ( );
FILL FILL_7_AND2X2_16 ( );
FILL FILL_8_AND2X2_16 ( );
FILL FILL_0_BUFX2_84 ( );
FILL FILL_1_BUFX2_84 ( );
FILL FILL_2_BUFX2_84 ( );
FILL FILL_3_BUFX2_84 ( );
FILL FILL_4_BUFX2_84 ( );
FILL FILL_5_BUFX2_84 ( );
FILL FILL_6_BUFX2_84 ( );
FILL FILL_0_NAND2X1_34 ( );
FILL FILL_1_NAND2X1_34 ( );
FILL FILL_2_NAND2X1_34 ( );
FILL FILL_3_NAND2X1_34 ( );
FILL FILL_4_NAND2X1_34 ( );
FILL FILL_5_NAND2X1_34 ( );
FILL FILL_6_NAND2X1_34 ( );
FILL FILL_0_NOR3X1_4 ( );
FILL FILL_1_NOR3X1_4 ( );
FILL FILL_2_NOR3X1_4 ( );
FILL FILL_3_NOR3X1_4 ( );
FILL FILL_4_NOR3X1_4 ( );
FILL FILL_5_NOR3X1_4 ( );
FILL FILL_6_NOR3X1_4 ( );
FILL FILL_7_NOR3X1_4 ( );
FILL FILL_8_NOR3X1_4 ( );
FILL FILL_9_NOR3X1_4 ( );
FILL FILL_10_NOR3X1_4 ( );
FILL FILL_11_NOR3X1_4 ( );
FILL FILL_12_NOR3X1_4 ( );
FILL FILL_13_NOR3X1_4 ( );
FILL FILL_14_NOR3X1_4 ( );
FILL FILL_15_NOR3X1_4 ( );
FILL FILL_16_NOR3X1_4 ( );
FILL FILL_17_NOR3X1_4 ( );
FILL FILL_18_NOR3X1_4 ( );
FILL FILL_0_DFFSR_114 ( );
FILL FILL_1_DFFSR_114 ( );
FILL FILL_2_DFFSR_114 ( );
FILL FILL_3_DFFSR_114 ( );
FILL FILL_4_DFFSR_114 ( );
FILL FILL_5_DFFSR_114 ( );
FILL FILL_6_DFFSR_114 ( );
FILL FILL_7_DFFSR_114 ( );
FILL FILL_8_DFFSR_114 ( );
FILL FILL_9_DFFSR_114 ( );
FILL FILL_10_DFFSR_114 ( );
FILL FILL_11_DFFSR_114 ( );
FILL FILL_12_DFFSR_114 ( );
FILL FILL_13_DFFSR_114 ( );
FILL FILL_14_DFFSR_114 ( );
FILL FILL_15_DFFSR_114 ( );
FILL FILL_16_DFFSR_114 ( );
FILL FILL_17_DFFSR_114 ( );
FILL FILL_18_DFFSR_114 ( );
FILL FILL_19_DFFSR_114 ( );
FILL FILL_20_DFFSR_114 ( );
FILL FILL_21_DFFSR_114 ( );
FILL FILL_22_DFFSR_114 ( );
FILL FILL_23_DFFSR_114 ( );
FILL FILL_24_DFFSR_114 ( );
FILL FILL_25_DFFSR_114 ( );
FILL FILL_26_DFFSR_114 ( );
FILL FILL_27_DFFSR_114 ( );
FILL FILL_28_DFFSR_114 ( );
FILL FILL_29_DFFSR_114 ( );
FILL FILL_30_DFFSR_114 ( );
FILL FILL_31_DFFSR_114 ( );
FILL FILL_32_DFFSR_114 ( );
FILL FILL_33_DFFSR_114 ( );
FILL FILL_34_DFFSR_114 ( );
FILL FILL_35_DFFSR_114 ( );
FILL FILL_36_DFFSR_114 ( );
FILL FILL_37_DFFSR_114 ( );
FILL FILL_38_DFFSR_114 ( );
FILL FILL_39_DFFSR_114 ( );
FILL FILL_40_DFFSR_114 ( );
FILL FILL_41_DFFSR_114 ( );
FILL FILL_42_DFFSR_114 ( );
FILL FILL_43_DFFSR_114 ( );
FILL FILL_44_DFFSR_114 ( );
FILL FILL_45_DFFSR_114 ( );
FILL FILL_46_DFFSR_114 ( );
FILL FILL_47_DFFSR_114 ( );
FILL FILL_48_DFFSR_114 ( );
FILL FILL_49_DFFSR_114 ( );
FILL FILL_50_DFFSR_114 ( );
FILL FILL_51_DFFSR_114 ( );
FILL FILL_0_BUFX2_33 ( );
FILL FILL_1_BUFX2_33 ( );
FILL FILL_2_BUFX2_33 ( );
FILL FILL_3_BUFX2_33 ( );
FILL FILL_4_BUFX2_33 ( );
FILL FILL_5_BUFX2_33 ( );
FILL FILL_6_BUFX2_33 ( );
FILL FILL_0_NAND3X1_80 ( );
FILL FILL_1_NAND3X1_80 ( );
FILL FILL_2_NAND3X1_80 ( );
FILL FILL_3_NAND3X1_80 ( );
FILL FILL_4_NAND3X1_80 ( );
FILL FILL_5_NAND3X1_80 ( );
FILL FILL_6_NAND3X1_80 ( );
FILL FILL_7_NAND3X1_80 ( );
FILL FILL_8_NAND3X1_80 ( );
FILL FILL_0_NOR2X1_40 ( );
FILL FILL_1_NOR2X1_40 ( );
FILL FILL_2_NOR2X1_40 ( );
FILL FILL_3_NOR2X1_40 ( );
FILL FILL_4_NOR2X1_40 ( );
FILL FILL_5_NOR2X1_40 ( );
FILL FILL_6_NOR2X1_40 ( );
FILL FILL_0_NAND3X1_79 ( );
FILL FILL_1_NAND3X1_79 ( );
FILL FILL_2_NAND3X1_79 ( );
FILL FILL_3_NAND3X1_79 ( );
FILL FILL_4_NAND3X1_79 ( );
FILL FILL_5_NAND3X1_79 ( );
FILL FILL_6_NAND3X1_79 ( );
FILL FILL_7_NAND3X1_79 ( );
FILL FILL_8_NAND3X1_79 ( );
FILL FILL_9_NAND3X1_79 ( );
FILL FILL_0_AOI22X1_10 ( );
FILL FILL_1_AOI22X1_10 ( );
FILL FILL_2_AOI22X1_10 ( );
FILL FILL_3_AOI22X1_10 ( );
FILL FILL_4_AOI22X1_10 ( );
FILL FILL_5_AOI22X1_10 ( );
FILL FILL_6_AOI22X1_10 ( );
FILL FILL_7_AOI22X1_10 ( );
FILL FILL_8_AOI22X1_10 ( );
FILL FILL_9_AOI22X1_10 ( );
FILL FILL_10_AOI22X1_10 ( );
FILL FILL_0_DFFSR_202 ( );
FILL FILL_1_DFFSR_202 ( );
FILL FILL_2_DFFSR_202 ( );
FILL FILL_3_DFFSR_202 ( );
FILL FILL_4_DFFSR_202 ( );
FILL FILL_5_DFFSR_202 ( );
FILL FILL_6_DFFSR_202 ( );
FILL FILL_7_DFFSR_202 ( );
FILL FILL_8_DFFSR_202 ( );
FILL FILL_9_DFFSR_202 ( );
FILL FILL_10_DFFSR_202 ( );
FILL FILL_11_DFFSR_202 ( );
FILL FILL_12_DFFSR_202 ( );
FILL FILL_13_DFFSR_202 ( );
FILL FILL_14_DFFSR_202 ( );
FILL FILL_15_DFFSR_202 ( );
FILL FILL_16_DFFSR_202 ( );
FILL FILL_17_DFFSR_202 ( );
FILL FILL_18_DFFSR_202 ( );
FILL FILL_19_DFFSR_202 ( );
FILL FILL_20_DFFSR_202 ( );
FILL FILL_21_DFFSR_202 ( );
FILL FILL_22_DFFSR_202 ( );
FILL FILL_23_DFFSR_202 ( );
FILL FILL_24_DFFSR_202 ( );
FILL FILL_25_DFFSR_202 ( );
FILL FILL_26_DFFSR_202 ( );
FILL FILL_27_DFFSR_202 ( );
FILL FILL_28_DFFSR_202 ( );
FILL FILL_29_DFFSR_202 ( );
FILL FILL_30_DFFSR_202 ( );
FILL FILL_31_DFFSR_202 ( );
FILL FILL_32_DFFSR_202 ( );
FILL FILL_33_DFFSR_202 ( );
FILL FILL_34_DFFSR_202 ( );
FILL FILL_35_DFFSR_202 ( );
FILL FILL_36_DFFSR_202 ( );
FILL FILL_37_DFFSR_202 ( );
FILL FILL_38_DFFSR_202 ( );
FILL FILL_39_DFFSR_202 ( );
FILL FILL_40_DFFSR_202 ( );
FILL FILL_41_DFFSR_202 ( );
FILL FILL_42_DFFSR_202 ( );
FILL FILL_43_DFFSR_202 ( );
FILL FILL_44_DFFSR_202 ( );
FILL FILL_45_DFFSR_202 ( );
FILL FILL_46_DFFSR_202 ( );
FILL FILL_47_DFFSR_202 ( );
FILL FILL_48_DFFSR_202 ( );
FILL FILL_49_DFFSR_202 ( );
FILL FILL_50_DFFSR_202 ( );
FILL FILL_51_DFFSR_202 ( );
FILL FILL_0_NAND2X1_95 ( );
FILL FILL_1_NAND2X1_95 ( );
FILL FILL_2_NAND2X1_95 ( );
FILL FILL_3_NAND2X1_95 ( );
FILL FILL_4_NAND2X1_95 ( );
FILL FILL_5_NAND2X1_95 ( );
FILL FILL_6_NAND2X1_95 ( );
FILL FILL_0_NAND2X1_109 ( );
FILL FILL_1_NAND2X1_109 ( );
FILL FILL_2_NAND2X1_109 ( );
FILL FILL_3_NAND2X1_109 ( );
FILL FILL_4_NAND2X1_109 ( );
FILL FILL_5_NAND2X1_109 ( );
FILL FILL_6_NAND2X1_109 ( );
FILL FILL_0_NAND2X1_93 ( );
FILL FILL_1_NAND2X1_93 ( );
FILL FILL_2_NAND2X1_93 ( );
FILL FILL_3_NAND2X1_93 ( );
FILL FILL_4_NAND2X1_93 ( );
FILL FILL_5_NAND2X1_93 ( );
FILL FILL_6_NAND2X1_93 ( );
FILL FILL_0_NAND3X1_173 ( );
FILL FILL_1_NAND3X1_173 ( );
FILL FILL_2_NAND3X1_173 ( );
FILL FILL_3_NAND3X1_173 ( );
FILL FILL_4_NAND3X1_173 ( );
FILL FILL_5_NAND3X1_173 ( );
FILL FILL_6_NAND3X1_173 ( );
FILL FILL_7_NAND3X1_173 ( );
FILL FILL_8_NAND3X1_173 ( );
FILL FILL_9_NAND3X1_173 ( );
FILL FILL_0_OAI21X1_66 ( );
FILL FILL_1_OAI21X1_66 ( );
FILL FILL_2_OAI21X1_66 ( );
FILL FILL_3_OAI21X1_66 ( );
FILL FILL_4_OAI21X1_66 ( );
FILL FILL_5_OAI21X1_66 ( );
FILL FILL_6_OAI21X1_66 ( );
FILL FILL_7_OAI21X1_66 ( );
FILL FILL_8_OAI21X1_66 ( );
FILL FILL_0_NOR2X1_70 ( );
FILL FILL_1_NOR2X1_70 ( );
FILL FILL_2_NOR2X1_70 ( );
FILL FILL_3_NOR2X1_70 ( );
FILL FILL_4_NOR2X1_70 ( );
FILL FILL_5_NOR2X1_70 ( );
FILL FILL_6_NOR2X1_70 ( );
FILL FILL_0_AND2X2_39 ( );
FILL FILL_1_AND2X2_39 ( );
FILL FILL_2_AND2X2_39 ( );
FILL FILL_3_AND2X2_39 ( );
FILL FILL_4_AND2X2_39 ( );
FILL FILL_5_AND2X2_39 ( );
FILL FILL_6_AND2X2_39 ( );
FILL FILL_7_AND2X2_39 ( );
FILL FILL_8_AND2X2_39 ( );
FILL FILL_0_DFFPOSX1_47 ( );
FILL FILL_1_DFFPOSX1_47 ( );
FILL FILL_2_DFFPOSX1_47 ( );
FILL FILL_3_DFFPOSX1_47 ( );
FILL FILL_4_DFFPOSX1_47 ( );
FILL FILL_5_DFFPOSX1_47 ( );
FILL FILL_6_DFFPOSX1_47 ( );
FILL FILL_7_DFFPOSX1_47 ( );
FILL FILL_8_DFFPOSX1_47 ( );
FILL FILL_9_DFFPOSX1_47 ( );
FILL FILL_10_DFFPOSX1_47 ( );
FILL FILL_11_DFFPOSX1_47 ( );
FILL FILL_12_DFFPOSX1_47 ( );
FILL FILL_13_DFFPOSX1_47 ( );
FILL FILL_14_DFFPOSX1_47 ( );
FILL FILL_15_DFFPOSX1_47 ( );
FILL FILL_16_DFFPOSX1_47 ( );
FILL FILL_17_DFFPOSX1_47 ( );
FILL FILL_18_DFFPOSX1_47 ( );
FILL FILL_19_DFFPOSX1_47 ( );
FILL FILL_20_DFFPOSX1_47 ( );
FILL FILL_21_DFFPOSX1_47 ( );
FILL FILL_22_DFFPOSX1_47 ( );
FILL FILL_23_DFFPOSX1_47 ( );
FILL FILL_24_DFFPOSX1_47 ( );
FILL FILL_25_DFFPOSX1_47 ( );
FILL FILL_26_DFFPOSX1_47 ( );
FILL FILL_27_DFFPOSX1_47 ( );
FILL FILL_0_INVX1_189 ( );
FILL FILL_1_INVX1_189 ( );
FILL FILL_2_INVX1_189 ( );
FILL FILL_3_INVX1_189 ( );
FILL FILL_4_INVX1_189 ( );
FILL FILL_0_NAND2X1_159 ( );
FILL FILL_1_NAND2X1_159 ( );
FILL FILL_2_NAND2X1_159 ( );
FILL FILL_3_NAND2X1_159 ( );
FILL FILL_4_NAND2X1_159 ( );
FILL FILL_5_NAND2X1_159 ( );
FILL FILL_6_NAND2X1_159 ( );
FILL FILL_0_DFFPOSX1_33 ( );
FILL FILL_1_DFFPOSX1_33 ( );
FILL FILL_2_DFFPOSX1_33 ( );
FILL FILL_3_DFFPOSX1_33 ( );
FILL FILL_4_DFFPOSX1_33 ( );
FILL FILL_5_DFFPOSX1_33 ( );
FILL FILL_6_DFFPOSX1_33 ( );
FILL FILL_7_DFFPOSX1_33 ( );
FILL FILL_8_DFFPOSX1_33 ( );
FILL FILL_9_DFFPOSX1_33 ( );
FILL FILL_10_DFFPOSX1_33 ( );
FILL FILL_11_DFFPOSX1_33 ( );
FILL FILL_12_DFFPOSX1_33 ( );
FILL FILL_13_DFFPOSX1_33 ( );
FILL FILL_14_DFFPOSX1_33 ( );
FILL FILL_15_DFFPOSX1_33 ( );
FILL FILL_16_DFFPOSX1_33 ( );
FILL FILL_17_DFFPOSX1_33 ( );
FILL FILL_18_DFFPOSX1_33 ( );
FILL FILL_19_DFFPOSX1_33 ( );
FILL FILL_20_DFFPOSX1_33 ( );
FILL FILL_21_DFFPOSX1_33 ( );
FILL FILL_22_DFFPOSX1_33 ( );
FILL FILL_23_DFFPOSX1_33 ( );
FILL FILL_24_DFFPOSX1_33 ( );
FILL FILL_25_DFFPOSX1_33 ( );
FILL FILL_26_DFFPOSX1_33 ( );
FILL FILL_27_DFFPOSX1_33 ( );
FILL FILL_0_DFFSR_71 ( );
FILL FILL_1_DFFSR_71 ( );
FILL FILL_2_DFFSR_71 ( );
FILL FILL_3_DFFSR_71 ( );
FILL FILL_4_DFFSR_71 ( );
FILL FILL_5_DFFSR_71 ( );
FILL FILL_6_DFFSR_71 ( );
FILL FILL_7_DFFSR_71 ( );
FILL FILL_8_DFFSR_71 ( );
FILL FILL_9_DFFSR_71 ( );
FILL FILL_10_DFFSR_71 ( );
FILL FILL_11_DFFSR_71 ( );
FILL FILL_12_DFFSR_71 ( );
FILL FILL_13_DFFSR_71 ( );
FILL FILL_14_DFFSR_71 ( );
FILL FILL_15_DFFSR_71 ( );
FILL FILL_16_DFFSR_71 ( );
FILL FILL_17_DFFSR_71 ( );
FILL FILL_18_DFFSR_71 ( );
FILL FILL_19_DFFSR_71 ( );
FILL FILL_20_DFFSR_71 ( );
FILL FILL_21_DFFSR_71 ( );
FILL FILL_22_DFFSR_71 ( );
FILL FILL_23_DFFSR_71 ( );
FILL FILL_24_DFFSR_71 ( );
FILL FILL_25_DFFSR_71 ( );
FILL FILL_26_DFFSR_71 ( );
FILL FILL_27_DFFSR_71 ( );
FILL FILL_28_DFFSR_71 ( );
FILL FILL_29_DFFSR_71 ( );
FILL FILL_30_DFFSR_71 ( );
FILL FILL_31_DFFSR_71 ( );
FILL FILL_32_DFFSR_71 ( );
FILL FILL_33_DFFSR_71 ( );
FILL FILL_34_DFFSR_71 ( );
FILL FILL_35_DFFSR_71 ( );
FILL FILL_36_DFFSR_71 ( );
FILL FILL_37_DFFSR_71 ( );
FILL FILL_38_DFFSR_71 ( );
FILL FILL_39_DFFSR_71 ( );
FILL FILL_40_DFFSR_71 ( );
FILL FILL_41_DFFSR_71 ( );
FILL FILL_42_DFFSR_71 ( );
FILL FILL_43_DFFSR_71 ( );
FILL FILL_44_DFFSR_71 ( );
FILL FILL_45_DFFSR_71 ( );
FILL FILL_46_DFFSR_71 ( );
FILL FILL_47_DFFSR_71 ( );
FILL FILL_48_DFFSR_71 ( );
FILL FILL_49_DFFSR_71 ( );
FILL FILL_50_DFFSR_71 ( );
FILL FILL_0_NAND2X1_174 ( );
FILL FILL_1_NAND2X1_174 ( );
FILL FILL_2_NAND2X1_174 ( );
FILL FILL_3_NAND2X1_174 ( );
FILL FILL_4_NAND2X1_174 ( );
FILL FILL_5_NAND2X1_174 ( );
FILL FILL_6_NAND2X1_174 ( );
FILL FILL_0_NAND2X1_175 ( );
FILL FILL_1_NAND2X1_175 ( );
FILL FILL_2_NAND2X1_175 ( );
FILL FILL_3_NAND2X1_175 ( );
FILL FILL_4_NAND2X1_175 ( );
FILL FILL_5_NAND2X1_175 ( );
FILL FILL_6_NAND2X1_175 ( );
FILL FILL_0_XOR2X1_11 ( );
FILL FILL_1_XOR2X1_11 ( );
FILL FILL_2_XOR2X1_11 ( );
FILL FILL_3_XOR2X1_11 ( );
FILL FILL_4_XOR2X1_11 ( );
FILL FILL_5_XOR2X1_11 ( );
FILL FILL_6_XOR2X1_11 ( );
FILL FILL_7_XOR2X1_11 ( );
FILL FILL_8_XOR2X1_11 ( );
FILL FILL_9_XOR2X1_11 ( );
FILL FILL_10_XOR2X1_11 ( );
FILL FILL_11_XOR2X1_11 ( );
FILL FILL_12_XOR2X1_11 ( );
FILL FILL_13_XOR2X1_11 ( );
FILL FILL_14_XOR2X1_11 ( );
FILL FILL_15_XOR2X1_11 ( );
FILL FILL_0_OAI21X1_116 ( );
FILL FILL_1_OAI21X1_116 ( );
FILL FILL_2_OAI21X1_116 ( );
FILL FILL_3_OAI21X1_116 ( );
FILL FILL_4_OAI21X1_116 ( );
FILL FILL_5_OAI21X1_116 ( );
FILL FILL_6_OAI21X1_116 ( );
FILL FILL_7_OAI21X1_116 ( );
FILL FILL_8_OAI21X1_116 ( );
FILL FILL_9_OAI21X1_116 ( );
FILL FILL_0_CLKBUF1_33 ( );
FILL FILL_1_CLKBUF1_33 ( );
FILL FILL_2_CLKBUF1_33 ( );
FILL FILL_3_CLKBUF1_33 ( );
FILL FILL_4_CLKBUF1_33 ( );
FILL FILL_5_CLKBUF1_33 ( );
FILL FILL_6_CLKBUF1_33 ( );
FILL FILL_7_CLKBUF1_33 ( );
FILL FILL_8_CLKBUF1_33 ( );
FILL FILL_9_CLKBUF1_33 ( );
FILL FILL_10_CLKBUF1_33 ( );
FILL FILL_11_CLKBUF1_33 ( );
FILL FILL_12_CLKBUF1_33 ( );
FILL FILL_13_CLKBUF1_33 ( );
FILL FILL_14_CLKBUF1_33 ( );
FILL FILL_15_CLKBUF1_33 ( );
FILL FILL_16_CLKBUF1_33 ( );
FILL FILL_17_CLKBUF1_33 ( );
FILL FILL_18_CLKBUF1_33 ( );
FILL FILL_19_CLKBUF1_33 ( );
FILL FILL_20_CLKBUF1_33 ( );
FILL FILL_0_DFFSR_91 ( );
FILL FILL_1_DFFSR_91 ( );
FILL FILL_2_DFFSR_91 ( );
FILL FILL_3_DFFSR_91 ( );
FILL FILL_4_DFFSR_91 ( );
FILL FILL_5_DFFSR_91 ( );
FILL FILL_6_DFFSR_91 ( );
FILL FILL_7_DFFSR_91 ( );
FILL FILL_8_DFFSR_91 ( );
FILL FILL_9_DFFSR_91 ( );
FILL FILL_10_DFFSR_91 ( );
FILL FILL_11_DFFSR_91 ( );
FILL FILL_12_DFFSR_91 ( );
FILL FILL_13_DFFSR_91 ( );
FILL FILL_14_DFFSR_91 ( );
FILL FILL_15_DFFSR_91 ( );
FILL FILL_16_DFFSR_91 ( );
FILL FILL_17_DFFSR_91 ( );
FILL FILL_18_DFFSR_91 ( );
FILL FILL_19_DFFSR_91 ( );
FILL FILL_20_DFFSR_91 ( );
FILL FILL_21_DFFSR_91 ( );
FILL FILL_22_DFFSR_91 ( );
FILL FILL_23_DFFSR_91 ( );
FILL FILL_24_DFFSR_91 ( );
FILL FILL_25_DFFSR_91 ( );
FILL FILL_26_DFFSR_91 ( );
FILL FILL_27_DFFSR_91 ( );
FILL FILL_28_DFFSR_91 ( );
FILL FILL_29_DFFSR_91 ( );
FILL FILL_30_DFFSR_91 ( );
FILL FILL_31_DFFSR_91 ( );
FILL FILL_32_DFFSR_91 ( );
FILL FILL_33_DFFSR_91 ( );
FILL FILL_34_DFFSR_91 ( );
FILL FILL_35_DFFSR_91 ( );
FILL FILL_36_DFFSR_91 ( );
FILL FILL_37_DFFSR_91 ( );
FILL FILL_38_DFFSR_91 ( );
FILL FILL_39_DFFSR_91 ( );
FILL FILL_40_DFFSR_91 ( );
FILL FILL_41_DFFSR_91 ( );
FILL FILL_42_DFFSR_91 ( );
FILL FILL_43_DFFSR_91 ( );
FILL FILL_44_DFFSR_91 ( );
FILL FILL_45_DFFSR_91 ( );
FILL FILL_46_DFFSR_91 ( );
FILL FILL_47_DFFSR_91 ( );
FILL FILL_48_DFFSR_91 ( );
FILL FILL_49_DFFSR_91 ( );
FILL FILL_50_DFFSR_91 ( );
FILL FILL_0_NOR2X1_3 ( );
FILL FILL_1_NOR2X1_3 ( );
FILL FILL_2_NOR2X1_3 ( );
FILL FILL_3_NOR2X1_3 ( );
FILL FILL_4_NOR2X1_3 ( );
FILL FILL_5_NOR2X1_3 ( );
FILL FILL_6_NOR2X1_3 ( );
FILL FILL_0_INVX1_63 ( );
FILL FILL_1_INVX1_63 ( );
FILL FILL_2_INVX1_63 ( );
FILL FILL_3_INVX1_63 ( );
FILL FILL_0_NAND2X1_33 ( );
FILL FILL_1_NAND2X1_33 ( );
FILL FILL_2_NAND2X1_33 ( );
FILL FILL_3_NAND2X1_33 ( );
FILL FILL_4_NAND2X1_33 ( );
FILL FILL_5_NAND2X1_33 ( );
FILL FILL_6_NAND2X1_33 ( );
FILL FILL_0_NOR2X1_34 ( );
FILL FILL_1_NOR2X1_34 ( );
FILL FILL_2_NOR2X1_34 ( );
FILL FILL_3_NOR2X1_34 ( );
FILL FILL_4_NOR2X1_34 ( );
FILL FILL_5_NOR2X1_34 ( );
FILL FILL_6_NOR2X1_34 ( );
FILL FILL_0_AND2X2_17 ( );
FILL FILL_1_AND2X2_17 ( );
FILL FILL_2_AND2X2_17 ( );
FILL FILL_3_AND2X2_17 ( );
FILL FILL_4_AND2X2_17 ( );
FILL FILL_5_AND2X2_17 ( );
FILL FILL_6_AND2X2_17 ( );
FILL FILL_7_AND2X2_17 ( );
FILL FILL_8_AND2X2_17 ( );
FILL FILL_0_DFFSR_106 ( );
FILL FILL_1_DFFSR_106 ( );
FILL FILL_2_DFFSR_106 ( );
FILL FILL_3_DFFSR_106 ( );
FILL FILL_4_DFFSR_106 ( );
FILL FILL_5_DFFSR_106 ( );
FILL FILL_6_DFFSR_106 ( );
FILL FILL_7_DFFSR_106 ( );
FILL FILL_8_DFFSR_106 ( );
FILL FILL_9_DFFSR_106 ( );
FILL FILL_10_DFFSR_106 ( );
FILL FILL_11_DFFSR_106 ( );
FILL FILL_12_DFFSR_106 ( );
FILL FILL_13_DFFSR_106 ( );
FILL FILL_14_DFFSR_106 ( );
FILL FILL_15_DFFSR_106 ( );
FILL FILL_16_DFFSR_106 ( );
FILL FILL_17_DFFSR_106 ( );
FILL FILL_18_DFFSR_106 ( );
FILL FILL_19_DFFSR_106 ( );
FILL FILL_20_DFFSR_106 ( );
FILL FILL_21_DFFSR_106 ( );
FILL FILL_22_DFFSR_106 ( );
FILL FILL_23_DFFSR_106 ( );
FILL FILL_24_DFFSR_106 ( );
FILL FILL_25_DFFSR_106 ( );
FILL FILL_26_DFFSR_106 ( );
FILL FILL_27_DFFSR_106 ( );
FILL FILL_28_DFFSR_106 ( );
FILL FILL_29_DFFSR_106 ( );
FILL FILL_30_DFFSR_106 ( );
FILL FILL_31_DFFSR_106 ( );
FILL FILL_32_DFFSR_106 ( );
FILL FILL_33_DFFSR_106 ( );
FILL FILL_34_DFFSR_106 ( );
FILL FILL_35_DFFSR_106 ( );
FILL FILL_36_DFFSR_106 ( );
FILL FILL_37_DFFSR_106 ( );
FILL FILL_38_DFFSR_106 ( );
FILL FILL_39_DFFSR_106 ( );
FILL FILL_40_DFFSR_106 ( );
FILL FILL_41_DFFSR_106 ( );
FILL FILL_42_DFFSR_106 ( );
FILL FILL_43_DFFSR_106 ( );
FILL FILL_44_DFFSR_106 ( );
FILL FILL_45_DFFSR_106 ( );
FILL FILL_46_DFFSR_106 ( );
FILL FILL_47_DFFSR_106 ( );
FILL FILL_48_DFFSR_106 ( );
FILL FILL_49_DFFSR_106 ( );
FILL FILL_50_DFFSR_106 ( );
FILL FILL_0_CLKBUF1_29 ( );
FILL FILL_1_CLKBUF1_29 ( );
FILL FILL_2_CLKBUF1_29 ( );
FILL FILL_3_CLKBUF1_29 ( );
FILL FILL_4_CLKBUF1_29 ( );
FILL FILL_5_CLKBUF1_29 ( );
FILL FILL_6_CLKBUF1_29 ( );
FILL FILL_7_CLKBUF1_29 ( );
FILL FILL_8_CLKBUF1_29 ( );
FILL FILL_9_CLKBUF1_29 ( );
FILL FILL_10_CLKBUF1_29 ( );
FILL FILL_11_CLKBUF1_29 ( );
FILL FILL_12_CLKBUF1_29 ( );
FILL FILL_13_CLKBUF1_29 ( );
FILL FILL_14_CLKBUF1_29 ( );
FILL FILL_15_CLKBUF1_29 ( );
FILL FILL_16_CLKBUF1_29 ( );
FILL FILL_17_CLKBUF1_29 ( );
FILL FILL_18_CLKBUF1_29 ( );
FILL FILL_19_CLKBUF1_29 ( );
FILL FILL_20_CLKBUF1_29 ( );
FILL FILL_0_NAND3X1_101 ( );
FILL FILL_1_NAND3X1_101 ( );
FILL FILL_2_NAND3X1_101 ( );
FILL FILL_3_NAND3X1_101 ( );
FILL FILL_4_NAND3X1_101 ( );
FILL FILL_5_NAND3X1_101 ( );
FILL FILL_6_NAND3X1_101 ( );
FILL FILL_7_NAND3X1_101 ( );
FILL FILL_8_NAND3X1_101 ( );
FILL FILL_0_NOR2X1_57 ( );
FILL FILL_1_NOR2X1_57 ( );
FILL FILL_2_NOR2X1_57 ( );
FILL FILL_3_NOR2X1_57 ( );
FILL FILL_4_NOR2X1_57 ( );
FILL FILL_5_NOR2X1_57 ( );
FILL FILL_6_NOR2X1_57 ( );
FILL FILL_0_OAI22X1_48 ( );
FILL FILL_1_OAI22X1_48 ( );
FILL FILL_2_OAI22X1_48 ( );
FILL FILL_3_OAI22X1_48 ( );
FILL FILL_4_OAI22X1_48 ( );
FILL FILL_5_OAI22X1_48 ( );
FILL FILL_6_OAI22X1_48 ( );
FILL FILL_7_OAI22X1_48 ( );
FILL FILL_8_OAI22X1_48 ( );
FILL FILL_9_OAI22X1_48 ( );
FILL FILL_10_OAI22X1_48 ( );
FILL FILL_0_INVX1_115 ( );
FILL FILL_1_INVX1_115 ( );
FILL FILL_2_INVX1_115 ( );
FILL FILL_3_INVX1_115 ( );
FILL FILL_4_INVX1_115 ( );
FILL FILL_0_DFFSR_141 ( );
FILL FILL_1_DFFSR_141 ( );
FILL FILL_2_DFFSR_141 ( );
FILL FILL_3_DFFSR_141 ( );
FILL FILL_4_DFFSR_141 ( );
FILL FILL_5_DFFSR_141 ( );
FILL FILL_6_DFFSR_141 ( );
FILL FILL_7_DFFSR_141 ( );
FILL FILL_8_DFFSR_141 ( );
FILL FILL_9_DFFSR_141 ( );
FILL FILL_10_DFFSR_141 ( );
FILL FILL_11_DFFSR_141 ( );
FILL FILL_12_DFFSR_141 ( );
FILL FILL_13_DFFSR_141 ( );
FILL FILL_14_DFFSR_141 ( );
FILL FILL_15_DFFSR_141 ( );
FILL FILL_16_DFFSR_141 ( );
FILL FILL_17_DFFSR_141 ( );
FILL FILL_18_DFFSR_141 ( );
FILL FILL_19_DFFSR_141 ( );
FILL FILL_20_DFFSR_141 ( );
FILL FILL_21_DFFSR_141 ( );
FILL FILL_22_DFFSR_141 ( );
FILL FILL_23_DFFSR_141 ( );
FILL FILL_24_DFFSR_141 ( );
FILL FILL_25_DFFSR_141 ( );
FILL FILL_26_DFFSR_141 ( );
FILL FILL_27_DFFSR_141 ( );
FILL FILL_28_DFFSR_141 ( );
FILL FILL_29_DFFSR_141 ( );
FILL FILL_30_DFFSR_141 ( );
FILL FILL_31_DFFSR_141 ( );
FILL FILL_32_DFFSR_141 ( );
FILL FILL_33_DFFSR_141 ( );
FILL FILL_34_DFFSR_141 ( );
FILL FILL_35_DFFSR_141 ( );
FILL FILL_36_DFFSR_141 ( );
FILL FILL_37_DFFSR_141 ( );
FILL FILL_38_DFFSR_141 ( );
FILL FILL_39_DFFSR_141 ( );
FILL FILL_40_DFFSR_141 ( );
FILL FILL_41_DFFSR_141 ( );
FILL FILL_42_DFFSR_141 ( );
FILL FILL_43_DFFSR_141 ( );
FILL FILL_44_DFFSR_141 ( );
FILL FILL_45_DFFSR_141 ( );
FILL FILL_46_DFFSR_141 ( );
FILL FILL_47_DFFSR_141 ( );
FILL FILL_48_DFFSR_141 ( );
FILL FILL_49_DFFSR_141 ( );
FILL FILL_50_DFFSR_141 ( );
FILL FILL_0_OAI21X1_63 ( );
FILL FILL_1_OAI21X1_63 ( );
FILL FILL_2_OAI21X1_63 ( );
FILL FILL_3_OAI21X1_63 ( );
FILL FILL_4_OAI21X1_63 ( );
FILL FILL_5_OAI21X1_63 ( );
FILL FILL_6_OAI21X1_63 ( );
FILL FILL_7_OAI21X1_63 ( );
FILL FILL_8_OAI21X1_63 ( );
FILL FILL_9_OAI21X1_63 ( );
FILL FILL_0_XOR2X1_4 ( );
FILL FILL_1_XOR2X1_4 ( );
FILL FILL_2_XOR2X1_4 ( );
FILL FILL_3_XOR2X1_4 ( );
FILL FILL_4_XOR2X1_4 ( );
FILL FILL_5_XOR2X1_4 ( );
FILL FILL_6_XOR2X1_4 ( );
FILL FILL_7_XOR2X1_4 ( );
FILL FILL_8_XOR2X1_4 ( );
FILL FILL_9_XOR2X1_4 ( );
FILL FILL_10_XOR2X1_4 ( );
FILL FILL_11_XOR2X1_4 ( );
FILL FILL_12_XOR2X1_4 ( );
FILL FILL_13_XOR2X1_4 ( );
FILL FILL_14_XOR2X1_4 ( );
FILL FILL_15_XOR2X1_4 ( );
FILL FILL_0_INVX1_160 ( );
FILL FILL_1_INVX1_160 ( );
FILL FILL_2_INVX1_160 ( );
FILL FILL_3_INVX1_160 ( );
FILL FILL_4_INVX1_160 ( );
FILL FILL_0_AOI21X1_30 ( );
FILL FILL_1_AOI21X1_30 ( );
FILL FILL_2_AOI21X1_30 ( );
FILL FILL_3_AOI21X1_30 ( );
FILL FILL_4_AOI21X1_30 ( );
FILL FILL_5_AOI21X1_30 ( );
FILL FILL_6_AOI21X1_30 ( );
FILL FILL_7_AOI21X1_30 ( );
FILL FILL_8_AOI21X1_30 ( );
FILL FILL_0_OAI21X1_50 ( );
FILL FILL_1_OAI21X1_50 ( );
FILL FILL_2_OAI21X1_50 ( );
FILL FILL_3_OAI21X1_50 ( );
FILL FILL_4_OAI21X1_50 ( );
FILL FILL_5_OAI21X1_50 ( );
FILL FILL_6_OAI21X1_50 ( );
FILL FILL_7_OAI21X1_50 ( );
FILL FILL_8_OAI21X1_50 ( );
FILL FILL_0_AND2X2_37 ( );
FILL FILL_1_AND2X2_37 ( );
FILL FILL_2_AND2X2_37 ( );
FILL FILL_3_AND2X2_37 ( );
FILL FILL_4_AND2X2_37 ( );
FILL FILL_5_AND2X2_37 ( );
FILL FILL_6_AND2X2_37 ( );
FILL FILL_7_AND2X2_37 ( );
FILL FILL_8_AND2X2_37 ( );
FILL FILL_0_AOI22X1_25 ( );
FILL FILL_1_AOI22X1_25 ( );
FILL FILL_2_AOI22X1_25 ( );
FILL FILL_3_AOI22X1_25 ( );
FILL FILL_4_AOI22X1_25 ( );
FILL FILL_5_AOI22X1_25 ( );
FILL FILL_6_AOI22X1_25 ( );
FILL FILL_7_AOI22X1_25 ( );
FILL FILL_8_AOI22X1_25 ( );
FILL FILL_9_AOI22X1_25 ( );
FILL FILL_10_AOI22X1_25 ( );
FILL FILL_11_AOI22X1_25 ( );
FILL FILL_0_DFFPOSX1_31 ( );
FILL FILL_1_DFFPOSX1_31 ( );
FILL FILL_2_DFFPOSX1_31 ( );
FILL FILL_3_DFFPOSX1_31 ( );
FILL FILL_4_DFFPOSX1_31 ( );
FILL FILL_5_DFFPOSX1_31 ( );
FILL FILL_6_DFFPOSX1_31 ( );
FILL FILL_7_DFFPOSX1_31 ( );
FILL FILL_8_DFFPOSX1_31 ( );
FILL FILL_9_DFFPOSX1_31 ( );
FILL FILL_10_DFFPOSX1_31 ( );
FILL FILL_11_DFFPOSX1_31 ( );
FILL FILL_12_DFFPOSX1_31 ( );
FILL FILL_13_DFFPOSX1_31 ( );
FILL FILL_14_DFFPOSX1_31 ( );
FILL FILL_15_DFFPOSX1_31 ( );
FILL FILL_16_DFFPOSX1_31 ( );
FILL FILL_17_DFFPOSX1_31 ( );
FILL FILL_18_DFFPOSX1_31 ( );
FILL FILL_19_DFFPOSX1_31 ( );
FILL FILL_20_DFFPOSX1_31 ( );
FILL FILL_21_DFFPOSX1_31 ( );
FILL FILL_22_DFFPOSX1_31 ( );
FILL FILL_23_DFFPOSX1_31 ( );
FILL FILL_24_DFFPOSX1_31 ( );
FILL FILL_25_DFFPOSX1_31 ( );
FILL FILL_26_DFFPOSX1_31 ( );
FILL FILL_27_DFFPOSX1_31 ( );
FILL FILL_0_NAND2X1_158 ( );
FILL FILL_1_NAND2X1_158 ( );
FILL FILL_2_NAND2X1_158 ( );
FILL FILL_3_NAND2X1_158 ( );
FILL FILL_4_NAND2X1_158 ( );
FILL FILL_5_NAND2X1_158 ( );
FILL FILL_6_NAND2X1_158 ( );
FILL FILL_0_AOI21X1_55 ( );
FILL FILL_1_AOI21X1_55 ( );
FILL FILL_2_AOI21X1_55 ( );
FILL FILL_3_AOI21X1_55 ( );
FILL FILL_4_AOI21X1_55 ( );
FILL FILL_5_AOI21X1_55 ( );
FILL FILL_6_AOI21X1_55 ( );
FILL FILL_7_AOI21X1_55 ( );
FILL FILL_8_AOI21X1_55 ( );
FILL FILL_0_DFFPOSX1_48 ( );
FILL FILL_1_DFFPOSX1_48 ( );
FILL FILL_2_DFFPOSX1_48 ( );
FILL FILL_3_DFFPOSX1_48 ( );
FILL FILL_4_DFFPOSX1_48 ( );
FILL FILL_5_DFFPOSX1_48 ( );
FILL FILL_6_DFFPOSX1_48 ( );
FILL FILL_7_DFFPOSX1_48 ( );
FILL FILL_8_DFFPOSX1_48 ( );
FILL FILL_9_DFFPOSX1_48 ( );
FILL FILL_10_DFFPOSX1_48 ( );
FILL FILL_11_DFFPOSX1_48 ( );
FILL FILL_12_DFFPOSX1_48 ( );
FILL FILL_13_DFFPOSX1_48 ( );
FILL FILL_14_DFFPOSX1_48 ( );
FILL FILL_15_DFFPOSX1_48 ( );
FILL FILL_16_DFFPOSX1_48 ( );
FILL FILL_17_DFFPOSX1_48 ( );
FILL FILL_18_DFFPOSX1_48 ( );
FILL FILL_19_DFFPOSX1_48 ( );
FILL FILL_20_DFFPOSX1_48 ( );
FILL FILL_21_DFFPOSX1_48 ( );
FILL FILL_22_DFFPOSX1_48 ( );
FILL FILL_23_DFFPOSX1_48 ( );
FILL FILL_24_DFFPOSX1_48 ( );
FILL FILL_25_DFFPOSX1_48 ( );
FILL FILL_26_DFFPOSX1_48 ( );
FILL FILL_27_DFFPOSX1_48 ( );
FILL FILL_0_AND2X2_4 ( );
FILL FILL_1_AND2X2_4 ( );
FILL FILL_2_AND2X2_4 ( );
FILL FILL_3_AND2X2_4 ( );
FILL FILL_4_AND2X2_4 ( );
FILL FILL_5_AND2X2_4 ( );
FILL FILL_6_AND2X2_4 ( );
FILL FILL_7_AND2X2_4 ( );
FILL FILL_8_AND2X2_4 ( );
FILL FILL_0_AND2X2_1 ( );
FILL FILL_1_AND2X2_1 ( );
FILL FILL_2_AND2X2_1 ( );
FILL FILL_3_AND2X2_1 ( );
FILL FILL_4_AND2X2_1 ( );
FILL FILL_5_AND2X2_1 ( );
FILL FILL_6_AND2X2_1 ( );
FILL FILL_7_AND2X2_1 ( );
FILL FILL_8_AND2X2_1 ( );
FILL FILL_9_AND2X2_1 ( );
FILL FILL_0_NOR2X1_82 ( );
FILL FILL_1_NOR2X1_82 ( );
FILL FILL_2_NOR2X1_82 ( );
FILL FILL_3_NOR2X1_82 ( );
FILL FILL_4_NOR2X1_82 ( );
FILL FILL_5_NOR2X1_82 ( );
FILL FILL_6_NOR2X1_82 ( );
FILL FILL_0_OAI21X1_117 ( );
FILL FILL_1_OAI21X1_117 ( );
FILL FILL_2_OAI21X1_117 ( );
FILL FILL_3_OAI21X1_117 ( );
FILL FILL_4_OAI21X1_117 ( );
FILL FILL_5_OAI21X1_117 ( );
FILL FILL_6_OAI21X1_117 ( );
FILL FILL_7_OAI21X1_117 ( );
FILL FILL_8_OAI21X1_117 ( );
FILL FILL_0_INVX1_214 ( );
FILL FILL_1_INVX1_214 ( );
FILL FILL_2_INVX1_214 ( );
FILL FILL_3_INVX1_214 ( );
FILL FILL_0_AOI21X1_68 ( );
FILL FILL_1_AOI21X1_68 ( );
FILL FILL_2_AOI21X1_68 ( );
FILL FILL_3_AOI21X1_68 ( );
FILL FILL_4_AOI21X1_68 ( );
FILL FILL_5_AOI21X1_68 ( );
FILL FILL_6_AOI21X1_68 ( );
FILL FILL_7_AOI21X1_68 ( );
FILL FILL_8_AOI21X1_68 ( );
FILL FILL_0_NAND2X1_176 ( );
FILL FILL_1_NAND2X1_176 ( );
FILL FILL_2_NAND2X1_176 ( );
FILL FILL_3_NAND2X1_176 ( );
FILL FILL_4_NAND2X1_176 ( );
FILL FILL_5_NAND2X1_176 ( );
FILL FILL_6_NAND2X1_176 ( );
FILL FILL_0_NAND2X1_177 ( );
FILL FILL_1_NAND2X1_177 ( );
FILL FILL_2_NAND2X1_177 ( );
FILL FILL_3_NAND2X1_177 ( );
FILL FILL_4_NAND2X1_177 ( );
FILL FILL_5_NAND2X1_177 ( );
FILL FILL_6_NAND2X1_177 ( );
FILL FILL_0_NOR2X1_81 ( );
FILL FILL_1_NOR2X1_81 ( );
FILL FILL_2_NOR2X1_81 ( );
FILL FILL_3_NOR2X1_81 ( );
FILL FILL_4_NOR2X1_81 ( );
FILL FILL_5_NOR2X1_81 ( );
FILL FILL_6_NOR2X1_81 ( );
FILL FILL_0_INVX1_217 ( );
FILL FILL_1_INVX1_217 ( );
FILL FILL_2_INVX1_217 ( );
FILL FILL_3_INVX1_217 ( );
FILL FILL_0_NOR2X1_12 ( );
FILL FILL_1_NOR2X1_12 ( );
FILL FILL_2_NOR2X1_12 ( );
FILL FILL_3_NOR2X1_12 ( );
FILL FILL_4_NOR2X1_12 ( );
FILL FILL_5_NOR2X1_12 ( );
FILL FILL_6_NOR2X1_12 ( );
FILL FILL_0_DFFSR_99 ( );
FILL FILL_1_DFFSR_99 ( );
FILL FILL_2_DFFSR_99 ( );
FILL FILL_3_DFFSR_99 ( );
FILL FILL_4_DFFSR_99 ( );
FILL FILL_5_DFFSR_99 ( );
FILL FILL_6_DFFSR_99 ( );
FILL FILL_7_DFFSR_99 ( );
FILL FILL_8_DFFSR_99 ( );
FILL FILL_9_DFFSR_99 ( );
FILL FILL_10_DFFSR_99 ( );
FILL FILL_11_DFFSR_99 ( );
FILL FILL_12_DFFSR_99 ( );
FILL FILL_13_DFFSR_99 ( );
FILL FILL_14_DFFSR_99 ( );
FILL FILL_15_DFFSR_99 ( );
FILL FILL_16_DFFSR_99 ( );
FILL FILL_17_DFFSR_99 ( );
FILL FILL_18_DFFSR_99 ( );
FILL FILL_19_DFFSR_99 ( );
FILL FILL_20_DFFSR_99 ( );
FILL FILL_21_DFFSR_99 ( );
FILL FILL_22_DFFSR_99 ( );
FILL FILL_23_DFFSR_99 ( );
FILL FILL_24_DFFSR_99 ( );
FILL FILL_25_DFFSR_99 ( );
FILL FILL_26_DFFSR_99 ( );
FILL FILL_27_DFFSR_99 ( );
FILL FILL_28_DFFSR_99 ( );
FILL FILL_29_DFFSR_99 ( );
FILL FILL_30_DFFSR_99 ( );
FILL FILL_31_DFFSR_99 ( );
FILL FILL_32_DFFSR_99 ( );
FILL FILL_33_DFFSR_99 ( );
FILL FILL_34_DFFSR_99 ( );
FILL FILL_35_DFFSR_99 ( );
FILL FILL_36_DFFSR_99 ( );
FILL FILL_37_DFFSR_99 ( );
FILL FILL_38_DFFSR_99 ( );
FILL FILL_39_DFFSR_99 ( );
FILL FILL_40_DFFSR_99 ( );
FILL FILL_41_DFFSR_99 ( );
FILL FILL_42_DFFSR_99 ( );
FILL FILL_43_DFFSR_99 ( );
FILL FILL_44_DFFSR_99 ( );
FILL FILL_45_DFFSR_99 ( );
FILL FILL_46_DFFSR_99 ( );
FILL FILL_47_DFFSR_99 ( );
FILL FILL_48_DFFSR_99 ( );
FILL FILL_49_DFFSR_99 ( );
FILL FILL_50_DFFSR_99 ( );
FILL FILL_0_BUFX2_85 ( );
FILL FILL_1_BUFX2_85 ( );
FILL FILL_2_BUFX2_85 ( );
FILL FILL_3_BUFX2_85 ( );
FILL FILL_4_BUFX2_85 ( );
FILL FILL_5_BUFX2_85 ( );
FILL FILL_6_BUFX2_85 ( );
FILL FILL_0_NAND3X1_8 ( );
FILL FILL_1_NAND3X1_8 ( );
FILL FILL_2_NAND3X1_8 ( );
FILL FILL_3_NAND3X1_8 ( );
FILL FILL_4_NAND3X1_8 ( );
FILL FILL_5_NAND3X1_8 ( );
FILL FILL_6_NAND3X1_8 ( );
FILL FILL_7_NAND3X1_8 ( );
FILL FILL_8_NAND3X1_8 ( );
FILL FILL_9_NAND3X1_8 ( );
FILL FILL_0_DFFSR_123 ( );
FILL FILL_1_DFFSR_123 ( );
FILL FILL_2_DFFSR_123 ( );
FILL FILL_3_DFFSR_123 ( );
FILL FILL_4_DFFSR_123 ( );
FILL FILL_5_DFFSR_123 ( );
FILL FILL_6_DFFSR_123 ( );
FILL FILL_7_DFFSR_123 ( );
FILL FILL_8_DFFSR_123 ( );
FILL FILL_9_DFFSR_123 ( );
FILL FILL_10_DFFSR_123 ( );
FILL FILL_11_DFFSR_123 ( );
FILL FILL_12_DFFSR_123 ( );
FILL FILL_13_DFFSR_123 ( );
FILL FILL_14_DFFSR_123 ( );
FILL FILL_15_DFFSR_123 ( );
FILL FILL_16_DFFSR_123 ( );
FILL FILL_17_DFFSR_123 ( );
FILL FILL_18_DFFSR_123 ( );
FILL FILL_19_DFFSR_123 ( );
FILL FILL_20_DFFSR_123 ( );
FILL FILL_21_DFFSR_123 ( );
FILL FILL_22_DFFSR_123 ( );
FILL FILL_23_DFFSR_123 ( );
FILL FILL_24_DFFSR_123 ( );
FILL FILL_25_DFFSR_123 ( );
FILL FILL_26_DFFSR_123 ( );
FILL FILL_27_DFFSR_123 ( );
FILL FILL_28_DFFSR_123 ( );
FILL FILL_29_DFFSR_123 ( );
FILL FILL_30_DFFSR_123 ( );
FILL FILL_31_DFFSR_123 ( );
FILL FILL_32_DFFSR_123 ( );
FILL FILL_33_DFFSR_123 ( );
FILL FILL_34_DFFSR_123 ( );
FILL FILL_35_DFFSR_123 ( );
FILL FILL_36_DFFSR_123 ( );
FILL FILL_37_DFFSR_123 ( );
FILL FILL_38_DFFSR_123 ( );
FILL FILL_39_DFFSR_123 ( );
FILL FILL_40_DFFSR_123 ( );
FILL FILL_41_DFFSR_123 ( );
FILL FILL_42_DFFSR_123 ( );
FILL FILL_43_DFFSR_123 ( );
FILL FILL_44_DFFSR_123 ( );
FILL FILL_45_DFFSR_123 ( );
FILL FILL_46_DFFSR_123 ( );
FILL FILL_47_DFFSR_123 ( );
FILL FILL_48_DFFSR_123 ( );
FILL FILL_49_DFFSR_123 ( );
FILL FILL_50_DFFSR_123 ( );
FILL FILL_51_DFFSR_123 ( );
FILL FILL_0_DFFSR_197 ( );
FILL FILL_1_DFFSR_197 ( );
FILL FILL_2_DFFSR_197 ( );
FILL FILL_3_DFFSR_197 ( );
FILL FILL_4_DFFSR_197 ( );
FILL FILL_5_DFFSR_197 ( );
FILL FILL_6_DFFSR_197 ( );
FILL FILL_7_DFFSR_197 ( );
FILL FILL_8_DFFSR_197 ( );
FILL FILL_9_DFFSR_197 ( );
FILL FILL_10_DFFSR_197 ( );
FILL FILL_11_DFFSR_197 ( );
FILL FILL_12_DFFSR_197 ( );
FILL FILL_13_DFFSR_197 ( );
FILL FILL_14_DFFSR_197 ( );
FILL FILL_15_DFFSR_197 ( );
FILL FILL_16_DFFSR_197 ( );
FILL FILL_17_DFFSR_197 ( );
FILL FILL_18_DFFSR_197 ( );
FILL FILL_19_DFFSR_197 ( );
FILL FILL_20_DFFSR_197 ( );
FILL FILL_21_DFFSR_197 ( );
FILL FILL_22_DFFSR_197 ( );
FILL FILL_23_DFFSR_197 ( );
FILL FILL_24_DFFSR_197 ( );
FILL FILL_25_DFFSR_197 ( );
FILL FILL_26_DFFSR_197 ( );
FILL FILL_27_DFFSR_197 ( );
FILL FILL_28_DFFSR_197 ( );
FILL FILL_29_DFFSR_197 ( );
FILL FILL_30_DFFSR_197 ( );
FILL FILL_31_DFFSR_197 ( );
FILL FILL_32_DFFSR_197 ( );
FILL FILL_33_DFFSR_197 ( );
FILL FILL_34_DFFSR_197 ( );
FILL FILL_35_DFFSR_197 ( );
FILL FILL_36_DFFSR_197 ( );
FILL FILL_37_DFFSR_197 ( );
FILL FILL_38_DFFSR_197 ( );
FILL FILL_39_DFFSR_197 ( );
FILL FILL_40_DFFSR_197 ( );
FILL FILL_41_DFFSR_197 ( );
FILL FILL_42_DFFSR_197 ( );
FILL FILL_43_DFFSR_197 ( );
FILL FILL_44_DFFSR_197 ( );
FILL FILL_45_DFFSR_197 ( );
FILL FILL_46_DFFSR_197 ( );
FILL FILL_47_DFFSR_197 ( );
FILL FILL_48_DFFSR_197 ( );
FILL FILL_49_DFFSR_197 ( );
FILL FILL_50_DFFSR_197 ( );
FILL FILL_0_NAND3X1_122 ( );
FILL FILL_1_NAND3X1_122 ( );
FILL FILL_2_NAND3X1_122 ( );
FILL FILL_3_NAND3X1_122 ( );
FILL FILL_4_NAND3X1_122 ( );
FILL FILL_5_NAND3X1_122 ( );
FILL FILL_6_NAND3X1_122 ( );
FILL FILL_7_NAND3X1_122 ( );
FILL FILL_8_NAND3X1_122 ( );
FILL FILL_0_NAND3X1_124 ( );
FILL FILL_1_NAND3X1_124 ( );
FILL FILL_2_NAND3X1_124 ( );
FILL FILL_3_NAND3X1_124 ( );
FILL FILL_4_NAND3X1_124 ( );
FILL FILL_5_NAND3X1_124 ( );
FILL FILL_6_NAND3X1_124 ( );
FILL FILL_7_NAND3X1_124 ( );
FILL FILL_8_NAND3X1_124 ( );
FILL FILL_0_OAI21X1_16 ( );
FILL FILL_1_OAI21X1_16 ( );
FILL FILL_2_OAI21X1_16 ( );
FILL FILL_3_OAI21X1_16 ( );
FILL FILL_4_OAI21X1_16 ( );
FILL FILL_5_OAI21X1_16 ( );
FILL FILL_6_OAI21X1_16 ( );
FILL FILL_7_OAI21X1_16 ( );
FILL FILL_8_OAI21X1_16 ( );
FILL FILL_0_NAND2X1_51 ( );
FILL FILL_1_NAND2X1_51 ( );
FILL FILL_2_NAND2X1_51 ( );
FILL FILL_3_NAND2X1_51 ( );
FILL FILL_4_NAND2X1_51 ( );
FILL FILL_5_NAND2X1_51 ( );
FILL FILL_6_NAND2X1_51 ( );
FILL FILL_0_DFFSR_160 ( );
FILL FILL_1_DFFSR_160 ( );
FILL FILL_2_DFFSR_160 ( );
FILL FILL_3_DFFSR_160 ( );
FILL FILL_4_DFFSR_160 ( );
FILL FILL_5_DFFSR_160 ( );
FILL FILL_6_DFFSR_160 ( );
FILL FILL_7_DFFSR_160 ( );
FILL FILL_8_DFFSR_160 ( );
FILL FILL_9_DFFSR_160 ( );
FILL FILL_10_DFFSR_160 ( );
FILL FILL_11_DFFSR_160 ( );
FILL FILL_12_DFFSR_160 ( );
FILL FILL_13_DFFSR_160 ( );
FILL FILL_14_DFFSR_160 ( );
FILL FILL_15_DFFSR_160 ( );
FILL FILL_16_DFFSR_160 ( );
FILL FILL_17_DFFSR_160 ( );
FILL FILL_18_DFFSR_160 ( );
FILL FILL_19_DFFSR_160 ( );
FILL FILL_20_DFFSR_160 ( );
FILL FILL_21_DFFSR_160 ( );
FILL FILL_22_DFFSR_160 ( );
FILL FILL_23_DFFSR_160 ( );
FILL FILL_24_DFFSR_160 ( );
FILL FILL_25_DFFSR_160 ( );
FILL FILL_26_DFFSR_160 ( );
FILL FILL_27_DFFSR_160 ( );
FILL FILL_28_DFFSR_160 ( );
FILL FILL_29_DFFSR_160 ( );
FILL FILL_30_DFFSR_160 ( );
FILL FILL_31_DFFSR_160 ( );
FILL FILL_32_DFFSR_160 ( );
FILL FILL_33_DFFSR_160 ( );
FILL FILL_34_DFFSR_160 ( );
FILL FILL_35_DFFSR_160 ( );
FILL FILL_36_DFFSR_160 ( );
FILL FILL_37_DFFSR_160 ( );
FILL FILL_38_DFFSR_160 ( );
FILL FILL_39_DFFSR_160 ( );
FILL FILL_40_DFFSR_160 ( );
FILL FILL_41_DFFSR_160 ( );
FILL FILL_42_DFFSR_160 ( );
FILL FILL_43_DFFSR_160 ( );
FILL FILL_44_DFFSR_160 ( );
FILL FILL_45_DFFSR_160 ( );
FILL FILL_46_DFFSR_160 ( );
FILL FILL_47_DFFSR_160 ( );
FILL FILL_48_DFFSR_160 ( );
FILL FILL_49_DFFSR_160 ( );
FILL FILL_50_DFFSR_160 ( );
FILL FILL_0_XNOR2X1_3 ( );
FILL FILL_1_XNOR2X1_3 ( );
FILL FILL_2_XNOR2X1_3 ( );
FILL FILL_3_XNOR2X1_3 ( );
FILL FILL_4_XNOR2X1_3 ( );
FILL FILL_5_XNOR2X1_3 ( );
FILL FILL_6_XNOR2X1_3 ( );
FILL FILL_7_XNOR2X1_3 ( );
FILL FILL_8_XNOR2X1_3 ( );
FILL FILL_9_XNOR2X1_3 ( );
FILL FILL_10_XNOR2X1_3 ( );
FILL FILL_11_XNOR2X1_3 ( );
FILL FILL_12_XNOR2X1_3 ( );
FILL FILL_13_XNOR2X1_3 ( );
FILL FILL_14_XNOR2X1_3 ( );
FILL FILL_15_XNOR2X1_3 ( );
FILL FILL_16_XNOR2X1_3 ( );
FILL FILL_0_AOI22X1_26 ( );
FILL FILL_1_AOI22X1_26 ( );
FILL FILL_2_AOI22X1_26 ( );
FILL FILL_3_AOI22X1_26 ( );
FILL FILL_4_AOI22X1_26 ( );
FILL FILL_5_AOI22X1_26 ( );
FILL FILL_6_AOI22X1_26 ( );
FILL FILL_7_AOI22X1_26 ( );
FILL FILL_8_AOI22X1_26 ( );
FILL FILL_9_AOI22X1_26 ( );
FILL FILL_10_AOI22X1_26 ( );
FILL FILL_11_AOI22X1_26 ( );
FILL FILL_0_NAND3X1_203 ( );
FILL FILL_1_NAND3X1_203 ( );
FILL FILL_2_NAND3X1_203 ( );
FILL FILL_3_NAND3X1_203 ( );
FILL FILL_4_NAND3X1_203 ( );
FILL FILL_5_NAND3X1_203 ( );
FILL FILL_6_NAND3X1_203 ( );
FILL FILL_7_NAND3X1_203 ( );
FILL FILL_8_NAND3X1_203 ( );
FILL FILL_0_NOR2X1_71 ( );
FILL FILL_1_NOR2X1_71 ( );
FILL FILL_2_NOR2X1_71 ( );
FILL FILL_3_NOR2X1_71 ( );
FILL FILL_4_NOR2X1_71 ( );
FILL FILL_5_NOR2X1_71 ( );
FILL FILL_6_NOR2X1_71 ( );
FILL FILL_0_OAI21X1_67 ( );
FILL FILL_1_OAI21X1_67 ( );
FILL FILL_2_OAI21X1_67 ( );
FILL FILL_3_OAI21X1_67 ( );
FILL FILL_4_OAI21X1_67 ( );
FILL FILL_5_OAI21X1_67 ( );
FILL FILL_6_OAI21X1_67 ( );
FILL FILL_7_OAI21X1_67 ( );
FILL FILL_8_OAI21X1_67 ( );
FILL FILL_0_NAND2X1_97 ( );
FILL FILL_1_NAND2X1_97 ( );
FILL FILL_2_NAND2X1_97 ( );
FILL FILL_3_NAND2X1_97 ( );
FILL FILL_4_NAND2X1_97 ( );
FILL FILL_5_NAND2X1_97 ( );
FILL FILL_6_NAND2X1_97 ( );
FILL FILL_0_NAND3X1_199 ( );
FILL FILL_1_NAND3X1_199 ( );
FILL FILL_2_NAND3X1_199 ( );
FILL FILL_3_NAND3X1_199 ( );
FILL FILL_4_NAND3X1_199 ( );
FILL FILL_5_NAND3X1_199 ( );
FILL FILL_6_NAND3X1_199 ( );
FILL FILL_7_NAND3X1_199 ( );
FILL FILL_8_NAND3X1_199 ( );
FILL FILL_0_BUFX2_40 ( );
FILL FILL_1_BUFX2_40 ( );
FILL FILL_2_BUFX2_40 ( );
FILL FILL_3_BUFX2_40 ( );
FILL FILL_4_BUFX2_40 ( );
FILL FILL_5_BUFX2_40 ( );
FILL FILL_6_BUFX2_40 ( );
FILL FILL_0_BUFX2_37 ( );
FILL FILL_1_BUFX2_37 ( );
FILL FILL_2_BUFX2_37 ( );
FILL FILL_3_BUFX2_37 ( );
FILL FILL_4_BUFX2_37 ( );
FILL FILL_5_BUFX2_37 ( );
FILL FILL_6_BUFX2_37 ( );
FILL FILL_0_NAND2X1_152 ( );
FILL FILL_1_NAND2X1_152 ( );
FILL FILL_2_NAND2X1_152 ( );
FILL FILL_3_NAND2X1_152 ( );
FILL FILL_4_NAND2X1_152 ( );
FILL FILL_5_NAND2X1_152 ( );
FILL FILL_6_NAND2X1_152 ( );
FILL FILL_0_NAND2X1_139 ( );
FILL FILL_1_NAND2X1_139 ( );
FILL FILL_2_NAND2X1_139 ( );
FILL FILL_3_NAND2X1_139 ( );
FILL FILL_4_NAND2X1_139 ( );
FILL FILL_5_NAND2X1_139 ( );
FILL FILL_6_NAND2X1_139 ( );
FILL FILL_0_DFFSR_100 ( );
FILL FILL_1_DFFSR_100 ( );
FILL FILL_2_DFFSR_100 ( );
FILL FILL_3_DFFSR_100 ( );
FILL FILL_4_DFFSR_100 ( );
FILL FILL_5_DFFSR_100 ( );
FILL FILL_6_DFFSR_100 ( );
FILL FILL_7_DFFSR_100 ( );
FILL FILL_8_DFFSR_100 ( );
FILL FILL_9_DFFSR_100 ( );
FILL FILL_10_DFFSR_100 ( );
FILL FILL_11_DFFSR_100 ( );
FILL FILL_12_DFFSR_100 ( );
FILL FILL_13_DFFSR_100 ( );
FILL FILL_14_DFFSR_100 ( );
FILL FILL_15_DFFSR_100 ( );
FILL FILL_16_DFFSR_100 ( );
FILL FILL_17_DFFSR_100 ( );
FILL FILL_18_DFFSR_100 ( );
FILL FILL_19_DFFSR_100 ( );
FILL FILL_20_DFFSR_100 ( );
FILL FILL_21_DFFSR_100 ( );
FILL FILL_22_DFFSR_100 ( );
FILL FILL_23_DFFSR_100 ( );
FILL FILL_24_DFFSR_100 ( );
FILL FILL_25_DFFSR_100 ( );
FILL FILL_26_DFFSR_100 ( );
FILL FILL_27_DFFSR_100 ( );
FILL FILL_28_DFFSR_100 ( );
FILL FILL_29_DFFSR_100 ( );
FILL FILL_30_DFFSR_100 ( );
FILL FILL_31_DFFSR_100 ( );
FILL FILL_32_DFFSR_100 ( );
FILL FILL_33_DFFSR_100 ( );
FILL FILL_34_DFFSR_100 ( );
FILL FILL_35_DFFSR_100 ( );
FILL FILL_36_DFFSR_100 ( );
FILL FILL_37_DFFSR_100 ( );
FILL FILL_38_DFFSR_100 ( );
FILL FILL_39_DFFSR_100 ( );
FILL FILL_40_DFFSR_100 ( );
FILL FILL_41_DFFSR_100 ( );
FILL FILL_42_DFFSR_100 ( );
FILL FILL_43_DFFSR_100 ( );
FILL FILL_44_DFFSR_100 ( );
FILL FILL_45_DFFSR_100 ( );
FILL FILL_46_DFFSR_100 ( );
FILL FILL_47_DFFSR_100 ( );
FILL FILL_48_DFFSR_100 ( );
FILL FILL_49_DFFSR_100 ( );
FILL FILL_50_DFFSR_100 ( );
FILL FILL_0_NOR2X1_2 ( );
FILL FILL_1_NOR2X1_2 ( );
FILL FILL_2_NOR2X1_2 ( );
FILL FILL_3_NOR2X1_2 ( );
FILL FILL_4_NOR2X1_2 ( );
FILL FILL_5_NOR2X1_2 ( );
FILL FILL_6_NOR2X1_2 ( );
FILL FILL_0_AOI21X1_69 ( );
FILL FILL_1_AOI21X1_69 ( );
FILL FILL_2_AOI21X1_69 ( );
FILL FILL_3_AOI21X1_69 ( );
FILL FILL_4_AOI21X1_69 ( );
FILL FILL_5_AOI21X1_69 ( );
FILL FILL_6_AOI21X1_69 ( );
FILL FILL_7_AOI21X1_69 ( );
FILL FILL_8_AOI21X1_69 ( );
FILL FILL_0_NAND2X1_179 ( );
FILL FILL_1_NAND2X1_179 ( );
FILL FILL_2_NAND2X1_179 ( );
FILL FILL_3_NAND2X1_179 ( );
FILL FILL_4_NAND2X1_179 ( );
FILL FILL_5_NAND2X1_179 ( );
FILL FILL_6_NAND2X1_179 ( );
FILL FILL_0_NAND2X1_180 ( );
FILL FILL_1_NAND2X1_180 ( );
FILL FILL_2_NAND2X1_180 ( );
FILL FILL_3_NAND2X1_180 ( );
FILL FILL_4_NAND2X1_180 ( );
FILL FILL_5_NAND2X1_180 ( );
FILL FILL_6_NAND2X1_180 ( );
FILL FILL_0_INVX1_212 ( );
FILL FILL_1_INVX1_212 ( );
FILL FILL_2_INVX1_212 ( );
FILL FILL_3_INVX1_212 ( );
FILL FILL_0_XOR2X1_13 ( );
FILL FILL_1_XOR2X1_13 ( );
FILL FILL_2_XOR2X1_13 ( );
FILL FILL_3_XOR2X1_13 ( );
FILL FILL_4_XOR2X1_13 ( );
FILL FILL_5_XOR2X1_13 ( );
FILL FILL_6_XOR2X1_13 ( );
FILL FILL_7_XOR2X1_13 ( );
FILL FILL_8_XOR2X1_13 ( );
FILL FILL_9_XOR2X1_13 ( );
FILL FILL_10_XOR2X1_13 ( );
FILL FILL_11_XOR2X1_13 ( );
FILL FILL_12_XOR2X1_13 ( );
FILL FILL_13_XOR2X1_13 ( );
FILL FILL_14_XOR2X1_13 ( );
FILL FILL_15_XOR2X1_13 ( );
FILL FILL_16_XOR2X1_13 ( );
FILL FILL_0_INVX1_216 ( );
FILL FILL_1_INVX1_216 ( );
FILL FILL_2_INVX1_216 ( );
FILL FILL_3_INVX1_216 ( );
FILL FILL_4_INVX1_216 ( );
FILL FILL_0_NOR2X1_14 ( );
FILL FILL_1_NOR2X1_14 ( );
FILL FILL_2_NOR2X1_14 ( );
FILL FILL_3_NOR2X1_14 ( );
FILL FILL_4_NOR2X1_14 ( );
FILL FILL_5_NOR2X1_14 ( );
FILL FILL_6_NOR2X1_14 ( );
FILL FILL_0_NAND3X1_24 ( );
FILL FILL_1_NAND3X1_24 ( );
FILL FILL_2_NAND3X1_24 ( );
FILL FILL_3_NAND3X1_24 ( );
FILL FILL_4_NAND3X1_24 ( );
FILL FILL_5_NAND3X1_24 ( );
FILL FILL_6_NAND3X1_24 ( );
FILL FILL_7_NAND3X1_24 ( );
FILL FILL_8_NAND3X1_24 ( );
FILL FILL_9_NAND3X1_24 ( );
FILL FILL_0_BUFX2_89 ( );
FILL FILL_1_BUFX2_89 ( );
FILL FILL_2_BUFX2_89 ( );
FILL FILL_3_BUFX2_89 ( );
FILL FILL_4_BUFX2_89 ( );
FILL FILL_5_BUFX2_89 ( );
FILL FILL_6_BUFX2_89 ( );
FILL FILL_0_AOI22X1_3 ( );
FILL FILL_1_AOI22X1_3 ( );
FILL FILL_2_AOI22X1_3 ( );
FILL FILL_3_AOI22X1_3 ( );
FILL FILL_4_AOI22X1_3 ( );
FILL FILL_5_AOI22X1_3 ( );
FILL FILL_6_AOI22X1_3 ( );
FILL FILL_7_AOI22X1_3 ( );
FILL FILL_8_AOI22X1_3 ( );
FILL FILL_9_AOI22X1_3 ( );
FILL FILL_10_AOI22X1_3 ( );
FILL FILL_11_AOI22X1_3 ( );
FILL FILL_0_DFFSR_97 ( );
FILL FILL_1_DFFSR_97 ( );
FILL FILL_2_DFFSR_97 ( );
FILL FILL_3_DFFSR_97 ( );
FILL FILL_4_DFFSR_97 ( );
FILL FILL_5_DFFSR_97 ( );
FILL FILL_6_DFFSR_97 ( );
FILL FILL_7_DFFSR_97 ( );
FILL FILL_8_DFFSR_97 ( );
FILL FILL_9_DFFSR_97 ( );
FILL FILL_10_DFFSR_97 ( );
FILL FILL_11_DFFSR_97 ( );
FILL FILL_12_DFFSR_97 ( );
FILL FILL_13_DFFSR_97 ( );
FILL FILL_14_DFFSR_97 ( );
FILL FILL_15_DFFSR_97 ( );
FILL FILL_16_DFFSR_97 ( );
FILL FILL_17_DFFSR_97 ( );
FILL FILL_18_DFFSR_97 ( );
FILL FILL_19_DFFSR_97 ( );
FILL FILL_20_DFFSR_97 ( );
FILL FILL_21_DFFSR_97 ( );
FILL FILL_22_DFFSR_97 ( );
FILL FILL_23_DFFSR_97 ( );
FILL FILL_24_DFFSR_97 ( );
FILL FILL_25_DFFSR_97 ( );
FILL FILL_26_DFFSR_97 ( );
FILL FILL_27_DFFSR_97 ( );
FILL FILL_28_DFFSR_97 ( );
FILL FILL_29_DFFSR_97 ( );
FILL FILL_30_DFFSR_97 ( );
FILL FILL_31_DFFSR_97 ( );
FILL FILL_32_DFFSR_97 ( );
FILL FILL_33_DFFSR_97 ( );
FILL FILL_34_DFFSR_97 ( );
FILL FILL_35_DFFSR_97 ( );
FILL FILL_36_DFFSR_97 ( );
FILL FILL_37_DFFSR_97 ( );
FILL FILL_38_DFFSR_97 ( );
FILL FILL_39_DFFSR_97 ( );
FILL FILL_40_DFFSR_97 ( );
FILL FILL_41_DFFSR_97 ( );
FILL FILL_42_DFFSR_97 ( );
FILL FILL_43_DFFSR_97 ( );
FILL FILL_44_DFFSR_97 ( );
FILL FILL_45_DFFSR_97 ( );
FILL FILL_46_DFFSR_97 ( );
FILL FILL_47_DFFSR_97 ( );
FILL FILL_48_DFFSR_97 ( );
FILL FILL_49_DFFSR_97 ( );
FILL FILL_50_DFFSR_97 ( );
FILL FILL_0_AOI22X1_1 ( );
FILL FILL_1_AOI22X1_1 ( );
FILL FILL_2_AOI22X1_1 ( );
FILL FILL_3_AOI22X1_1 ( );
FILL FILL_4_AOI22X1_1 ( );
FILL FILL_5_AOI22X1_1 ( );
FILL FILL_6_AOI22X1_1 ( );
FILL FILL_7_AOI22X1_1 ( );
FILL FILL_8_AOI22X1_1 ( );
FILL FILL_9_AOI22X1_1 ( );
FILL FILL_10_AOI22X1_1 ( );
FILL FILL_11_AOI22X1_1 ( );
FILL FILL_0_DFFSR_115 ( );
FILL FILL_1_DFFSR_115 ( );
FILL FILL_2_DFFSR_115 ( );
FILL FILL_3_DFFSR_115 ( );
FILL FILL_4_DFFSR_115 ( );
FILL FILL_5_DFFSR_115 ( );
FILL FILL_6_DFFSR_115 ( );
FILL FILL_7_DFFSR_115 ( );
FILL FILL_8_DFFSR_115 ( );
FILL FILL_9_DFFSR_115 ( );
FILL FILL_10_DFFSR_115 ( );
FILL FILL_11_DFFSR_115 ( );
FILL FILL_12_DFFSR_115 ( );
FILL FILL_13_DFFSR_115 ( );
FILL FILL_14_DFFSR_115 ( );
FILL FILL_15_DFFSR_115 ( );
FILL FILL_16_DFFSR_115 ( );
FILL FILL_17_DFFSR_115 ( );
FILL FILL_18_DFFSR_115 ( );
FILL FILL_19_DFFSR_115 ( );
FILL FILL_20_DFFSR_115 ( );
FILL FILL_21_DFFSR_115 ( );
FILL FILL_22_DFFSR_115 ( );
FILL FILL_23_DFFSR_115 ( );
FILL FILL_24_DFFSR_115 ( );
FILL FILL_25_DFFSR_115 ( );
FILL FILL_26_DFFSR_115 ( );
FILL FILL_27_DFFSR_115 ( );
FILL FILL_28_DFFSR_115 ( );
FILL FILL_29_DFFSR_115 ( );
FILL FILL_30_DFFSR_115 ( );
FILL FILL_31_DFFSR_115 ( );
FILL FILL_32_DFFSR_115 ( );
FILL FILL_33_DFFSR_115 ( );
FILL FILL_34_DFFSR_115 ( );
FILL FILL_35_DFFSR_115 ( );
FILL FILL_36_DFFSR_115 ( );
FILL FILL_37_DFFSR_115 ( );
FILL FILL_38_DFFSR_115 ( );
FILL FILL_39_DFFSR_115 ( );
FILL FILL_40_DFFSR_115 ( );
FILL FILL_41_DFFSR_115 ( );
FILL FILL_42_DFFSR_115 ( );
FILL FILL_43_DFFSR_115 ( );
FILL FILL_44_DFFSR_115 ( );
FILL FILL_45_DFFSR_115 ( );
FILL FILL_46_DFFSR_115 ( );
FILL FILL_47_DFFSR_115 ( );
FILL FILL_48_DFFSR_115 ( );
FILL FILL_49_DFFSR_115 ( );
FILL FILL_50_DFFSR_115 ( );
FILL FILL_0_BUFX2_49 ( );
FILL FILL_1_BUFX2_49 ( );
FILL FILL_2_BUFX2_49 ( );
FILL FILL_3_BUFX2_49 ( );
FILL FILL_4_BUFX2_49 ( );
FILL FILL_5_BUFX2_49 ( );
FILL FILL_6_BUFX2_49 ( );
FILL FILL_0_BUFX2_82 ( );
FILL FILL_1_BUFX2_82 ( );
FILL FILL_2_BUFX2_82 ( );
FILL FILL_3_BUFX2_82 ( );
FILL FILL_4_BUFX2_82 ( );
FILL FILL_5_BUFX2_82 ( );
FILL FILL_6_BUFX2_82 ( );
FILL FILL_0_CLKBUF1_27 ( );
FILL FILL_1_CLKBUF1_27 ( );
FILL FILL_2_CLKBUF1_27 ( );
FILL FILL_3_CLKBUF1_27 ( );
FILL FILL_4_CLKBUF1_27 ( );
FILL FILL_5_CLKBUF1_27 ( );
FILL FILL_6_CLKBUF1_27 ( );
FILL FILL_7_CLKBUF1_27 ( );
FILL FILL_8_CLKBUF1_27 ( );
FILL FILL_9_CLKBUF1_27 ( );
FILL FILL_10_CLKBUF1_27 ( );
FILL FILL_11_CLKBUF1_27 ( );
FILL FILL_12_CLKBUF1_27 ( );
FILL FILL_13_CLKBUF1_27 ( );
FILL FILL_14_CLKBUF1_27 ( );
FILL FILL_15_CLKBUF1_27 ( );
FILL FILL_16_CLKBUF1_27 ( );
FILL FILL_17_CLKBUF1_27 ( );
FILL FILL_18_CLKBUF1_27 ( );
FILL FILL_19_CLKBUF1_27 ( );
FILL FILL_20_CLKBUF1_27 ( );
FILL FILL_0_AND2X2_26 ( );
FILL FILL_1_AND2X2_26 ( );
FILL FILL_2_AND2X2_26 ( );
FILL FILL_3_AND2X2_26 ( );
FILL FILL_4_AND2X2_26 ( );
FILL FILL_5_AND2X2_26 ( );
FILL FILL_6_AND2X2_26 ( );
FILL FILL_7_AND2X2_26 ( );
FILL FILL_8_AND2X2_26 ( );
FILL FILL_9_AND2X2_26 ( );
FILL FILL_0_NAND3X1_74 ( );
FILL FILL_1_NAND3X1_74 ( );
FILL FILL_2_NAND3X1_74 ( );
FILL FILL_3_NAND3X1_74 ( );
FILL FILL_4_NAND3X1_74 ( );
FILL FILL_5_NAND3X1_74 ( );
FILL FILL_6_NAND3X1_74 ( );
FILL FILL_7_NAND3X1_74 ( );
FILL FILL_8_NAND3X1_74 ( );
FILL FILL_0_NAND3X1_73 ( );
FILL FILL_1_NAND3X1_73 ( );
FILL FILL_2_NAND3X1_73 ( );
FILL FILL_3_NAND3X1_73 ( );
FILL FILL_4_NAND3X1_73 ( );
FILL FILL_5_NAND3X1_73 ( );
FILL FILL_6_NAND3X1_73 ( );
FILL FILL_7_NAND3X1_73 ( );
FILL FILL_8_NAND3X1_73 ( );
FILL FILL_9_NAND3X1_73 ( );
FILL FILL_0_NAND3X1_121 ( );
FILL FILL_1_NAND3X1_121 ( );
FILL FILL_2_NAND3X1_121 ( );
FILL FILL_3_NAND3X1_121 ( );
FILL FILL_4_NAND3X1_121 ( );
FILL FILL_5_NAND3X1_121 ( );
FILL FILL_6_NAND3X1_121 ( );
FILL FILL_7_NAND3X1_121 ( );
FILL FILL_8_NAND3X1_121 ( );
FILL FILL_9_NAND3X1_121 ( );
FILL FILL_0_DFFSR_192 ( );
FILL FILL_1_DFFSR_192 ( );
FILL FILL_2_DFFSR_192 ( );
FILL FILL_3_DFFSR_192 ( );
FILL FILL_4_DFFSR_192 ( );
FILL FILL_5_DFFSR_192 ( );
FILL FILL_6_DFFSR_192 ( );
FILL FILL_7_DFFSR_192 ( );
FILL FILL_8_DFFSR_192 ( );
FILL FILL_9_DFFSR_192 ( );
FILL FILL_10_DFFSR_192 ( );
FILL FILL_11_DFFSR_192 ( );
FILL FILL_12_DFFSR_192 ( );
FILL FILL_13_DFFSR_192 ( );
FILL FILL_14_DFFSR_192 ( );
FILL FILL_15_DFFSR_192 ( );
FILL FILL_16_DFFSR_192 ( );
FILL FILL_17_DFFSR_192 ( );
FILL FILL_18_DFFSR_192 ( );
FILL FILL_19_DFFSR_192 ( );
FILL FILL_20_DFFSR_192 ( );
FILL FILL_21_DFFSR_192 ( );
FILL FILL_22_DFFSR_192 ( );
FILL FILL_23_DFFSR_192 ( );
FILL FILL_24_DFFSR_192 ( );
FILL FILL_25_DFFSR_192 ( );
FILL FILL_26_DFFSR_192 ( );
FILL FILL_27_DFFSR_192 ( );
FILL FILL_28_DFFSR_192 ( );
FILL FILL_29_DFFSR_192 ( );
FILL FILL_30_DFFSR_192 ( );
FILL FILL_31_DFFSR_192 ( );
FILL FILL_32_DFFSR_192 ( );
FILL FILL_33_DFFSR_192 ( );
FILL FILL_34_DFFSR_192 ( );
FILL FILL_35_DFFSR_192 ( );
FILL FILL_36_DFFSR_192 ( );
FILL FILL_37_DFFSR_192 ( );
FILL FILL_38_DFFSR_192 ( );
FILL FILL_39_DFFSR_192 ( );
FILL FILL_40_DFFSR_192 ( );
FILL FILL_41_DFFSR_192 ( );
FILL FILL_42_DFFSR_192 ( );
FILL FILL_43_DFFSR_192 ( );
FILL FILL_44_DFFSR_192 ( );
FILL FILL_45_DFFSR_192 ( );
FILL FILL_46_DFFSR_192 ( );
FILL FILL_47_DFFSR_192 ( );
FILL FILL_48_DFFSR_192 ( );
FILL FILL_49_DFFSR_192 ( );
FILL FILL_50_DFFSR_192 ( );
FILL FILL_0_OAI21X1_76 ( );
FILL FILL_1_OAI21X1_76 ( );
FILL FILL_2_OAI21X1_76 ( );
FILL FILL_3_OAI21X1_76 ( );
FILL FILL_4_OAI21X1_76 ( );
FILL FILL_5_OAI21X1_76 ( );
FILL FILL_6_OAI21X1_76 ( );
FILL FILL_7_OAI21X1_76 ( );
FILL FILL_8_OAI21X1_76 ( );
FILL FILL_0_OAI21X1_64 ( );
FILL FILL_1_OAI21X1_64 ( );
FILL FILL_2_OAI21X1_64 ( );
FILL FILL_3_OAI21X1_64 ( );
FILL FILL_4_OAI21X1_64 ( );
FILL FILL_5_OAI21X1_64 ( );
FILL FILL_6_OAI21X1_64 ( );
FILL FILL_7_OAI21X1_64 ( );
FILL FILL_8_OAI21X1_64 ( );
FILL FILL_0_AOI22X1_29 ( );
FILL FILL_1_AOI22X1_29 ( );
FILL FILL_2_AOI22X1_29 ( );
FILL FILL_3_AOI22X1_29 ( );
FILL FILL_4_AOI22X1_29 ( );
FILL FILL_5_AOI22X1_29 ( );
FILL FILL_6_AOI22X1_29 ( );
FILL FILL_7_AOI22X1_29 ( );
FILL FILL_8_AOI22X1_29 ( );
FILL FILL_9_AOI22X1_29 ( );
FILL FILL_10_AOI22X1_29 ( );
FILL FILL_11_AOI22X1_29 ( );
FILL FILL_0_NAND3X1_201 ( );
FILL FILL_1_NAND3X1_201 ( );
FILL FILL_2_NAND3X1_201 ( );
FILL FILL_3_NAND3X1_201 ( );
FILL FILL_4_NAND3X1_201 ( );
FILL FILL_5_NAND3X1_201 ( );
FILL FILL_6_NAND3X1_201 ( );
FILL FILL_7_NAND3X1_201 ( );
FILL FILL_8_NAND3X1_201 ( );
FILL FILL_9_NAND3X1_201 ( );
FILL FILL_0_NAND3X1_205 ( );
FILL FILL_1_NAND3X1_205 ( );
FILL FILL_2_NAND3X1_205 ( );
FILL FILL_3_NAND3X1_205 ( );
FILL FILL_4_NAND3X1_205 ( );
FILL FILL_5_NAND3X1_205 ( );
FILL FILL_6_NAND3X1_205 ( );
FILL FILL_7_NAND3X1_205 ( );
FILL FILL_8_NAND3X1_205 ( );
FILL FILL_0_INVX1_161 ( );
FILL FILL_1_INVX1_161 ( );
FILL FILL_2_INVX1_161 ( );
FILL FILL_3_INVX1_161 ( );
FILL FILL_4_INVX1_161 ( );
FILL FILL_0_OAI21X1_65 ( );
FILL FILL_1_OAI21X1_65 ( );
FILL FILL_2_OAI21X1_65 ( );
FILL FILL_3_OAI21X1_65 ( );
FILL FILL_4_OAI21X1_65 ( );
FILL FILL_5_OAI21X1_65 ( );
FILL FILL_6_OAI21X1_65 ( );
FILL FILL_7_OAI21X1_65 ( );
FILL FILL_8_OAI21X1_65 ( );
FILL FILL_0_DFFPOSX1_50 ( );
FILL FILL_1_DFFPOSX1_50 ( );
FILL FILL_2_DFFPOSX1_50 ( );
FILL FILL_3_DFFPOSX1_50 ( );
FILL FILL_4_DFFPOSX1_50 ( );
FILL FILL_5_DFFPOSX1_50 ( );
FILL FILL_6_DFFPOSX1_50 ( );
FILL FILL_7_DFFPOSX1_50 ( );
FILL FILL_8_DFFPOSX1_50 ( );
FILL FILL_9_DFFPOSX1_50 ( );
FILL FILL_10_DFFPOSX1_50 ( );
FILL FILL_11_DFFPOSX1_50 ( );
FILL FILL_12_DFFPOSX1_50 ( );
FILL FILL_13_DFFPOSX1_50 ( );
FILL FILL_14_DFFPOSX1_50 ( );
FILL FILL_15_DFFPOSX1_50 ( );
FILL FILL_16_DFFPOSX1_50 ( );
FILL FILL_17_DFFPOSX1_50 ( );
FILL FILL_18_DFFPOSX1_50 ( );
FILL FILL_19_DFFPOSX1_50 ( );
FILL FILL_20_DFFPOSX1_50 ( );
FILL FILL_21_DFFPOSX1_50 ( );
FILL FILL_22_DFFPOSX1_50 ( );
FILL FILL_23_DFFPOSX1_50 ( );
FILL FILL_24_DFFPOSX1_50 ( );
FILL FILL_25_DFFPOSX1_50 ( );
FILL FILL_26_DFFPOSX1_50 ( );
FILL FILL_27_DFFPOSX1_50 ( );
FILL FILL_0_NAND2X1_169 ( );
FILL FILL_1_NAND2X1_169 ( );
FILL FILL_2_NAND2X1_169 ( );
FILL FILL_3_NAND2X1_169 ( );
FILL FILL_4_NAND2X1_169 ( );
FILL FILL_5_NAND2X1_169 ( );
FILL FILL_6_NAND2X1_169 ( );
FILL FILL_0_OAI21X1_108 ( );
FILL FILL_1_OAI21X1_108 ( );
FILL FILL_2_OAI21X1_108 ( );
FILL FILL_3_OAI21X1_108 ( );
FILL FILL_4_OAI21X1_108 ( );
FILL FILL_5_OAI21X1_108 ( );
FILL FILL_6_OAI21X1_108 ( );
FILL FILL_7_OAI21X1_108 ( );
FILL FILL_8_OAI21X1_108 ( );
FILL FILL_0_INVX1_206 ( );
FILL FILL_1_INVX1_206 ( );
FILL FILL_2_INVX1_206 ( );
FILL FILL_3_INVX1_206 ( );
FILL FILL_4_INVX1_206 ( );
FILL FILL_0_NOR3X1_2 ( );
FILL FILL_1_NOR3X1_2 ( );
FILL FILL_2_NOR3X1_2 ( );
FILL FILL_3_NOR3X1_2 ( );
FILL FILL_4_NOR3X1_2 ( );
FILL FILL_5_NOR3X1_2 ( );
FILL FILL_6_NOR3X1_2 ( );
FILL FILL_7_NOR3X1_2 ( );
FILL FILL_8_NOR3X1_2 ( );
FILL FILL_9_NOR3X1_2 ( );
FILL FILL_10_NOR3X1_2 ( );
FILL FILL_11_NOR3X1_2 ( );
FILL FILL_12_NOR3X1_2 ( );
FILL FILL_13_NOR3X1_2 ( );
FILL FILL_14_NOR3X1_2 ( );
FILL FILL_15_NOR3X1_2 ( );
FILL FILL_16_NOR3X1_2 ( );
FILL FILL_17_NOR3X1_2 ( );
FILL FILL_0_NAND2X1_8 ( );
FILL FILL_1_NAND2X1_8 ( );
FILL FILL_2_NAND2X1_8 ( );
FILL FILL_3_NAND2X1_8 ( );
FILL FILL_4_NAND2X1_8 ( );
FILL FILL_5_NAND2X1_8 ( );
FILL FILL_6_NAND2X1_8 ( );
FILL FILL_0_NOR2X1_4 ( );
FILL FILL_1_NOR2X1_4 ( );
FILL FILL_2_NOR2X1_4 ( );
FILL FILL_3_NOR2X1_4 ( );
FILL FILL_4_NOR2X1_4 ( );
FILL FILL_5_NOR2X1_4 ( );
FILL FILL_6_NOR2X1_4 ( );
FILL FILL_0_AND2X2_3 ( );
FILL FILL_1_AND2X2_3 ( );
FILL FILL_2_AND2X2_3 ( );
FILL FILL_3_AND2X2_3 ( );
FILL FILL_4_AND2X2_3 ( );
FILL FILL_5_AND2X2_3 ( );
FILL FILL_6_AND2X2_3 ( );
FILL FILL_7_AND2X2_3 ( );
FILL FILL_8_AND2X2_3 ( );
FILL FILL_0_XOR2X1_14 ( );
FILL FILL_1_XOR2X1_14 ( );
FILL FILL_2_XOR2X1_14 ( );
FILL FILL_3_XOR2X1_14 ( );
FILL FILL_4_XOR2X1_14 ( );
FILL FILL_5_XOR2X1_14 ( );
FILL FILL_6_XOR2X1_14 ( );
FILL FILL_7_XOR2X1_14 ( );
FILL FILL_8_XOR2X1_14 ( );
FILL FILL_9_XOR2X1_14 ( );
FILL FILL_10_XOR2X1_14 ( );
FILL FILL_11_XOR2X1_14 ( );
FILL FILL_12_XOR2X1_14 ( );
FILL FILL_13_XOR2X1_14 ( );
FILL FILL_14_XOR2X1_14 ( );
FILL FILL_15_XOR2X1_14 ( );
FILL FILL_16_XOR2X1_14 ( );
FILL FILL_0_NAND2X1_178 ( );
FILL FILL_1_NAND2X1_178 ( );
FILL FILL_2_NAND2X1_178 ( );
FILL FILL_3_NAND2X1_178 ( );
FILL FILL_4_NAND2X1_178 ( );
FILL FILL_5_NAND2X1_178 ( );
FILL FILL_6_NAND2X1_178 ( );
FILL FILL_0_INVX1_30 ( );
FILL FILL_1_INVX1_30 ( );
FILL FILL_2_INVX1_30 ( );
FILL FILL_3_INVX1_30 ( );
FILL FILL_0_DFFSR_14 ( );
FILL FILL_1_DFFSR_14 ( );
FILL FILL_2_DFFSR_14 ( );
FILL FILL_3_DFFSR_14 ( );
FILL FILL_4_DFFSR_14 ( );
FILL FILL_5_DFFSR_14 ( );
FILL FILL_6_DFFSR_14 ( );
FILL FILL_7_DFFSR_14 ( );
FILL FILL_8_DFFSR_14 ( );
FILL FILL_9_DFFSR_14 ( );
FILL FILL_10_DFFSR_14 ( );
FILL FILL_11_DFFSR_14 ( );
FILL FILL_12_DFFSR_14 ( );
FILL FILL_13_DFFSR_14 ( );
FILL FILL_14_DFFSR_14 ( );
FILL FILL_15_DFFSR_14 ( );
FILL FILL_16_DFFSR_14 ( );
FILL FILL_17_DFFSR_14 ( );
FILL FILL_18_DFFSR_14 ( );
FILL FILL_19_DFFSR_14 ( );
FILL FILL_20_DFFSR_14 ( );
FILL FILL_21_DFFSR_14 ( );
FILL FILL_22_DFFSR_14 ( );
FILL FILL_23_DFFSR_14 ( );
FILL FILL_24_DFFSR_14 ( );
FILL FILL_25_DFFSR_14 ( );
FILL FILL_26_DFFSR_14 ( );
FILL FILL_27_DFFSR_14 ( );
FILL FILL_28_DFFSR_14 ( );
FILL FILL_29_DFFSR_14 ( );
FILL FILL_30_DFFSR_14 ( );
FILL FILL_31_DFFSR_14 ( );
FILL FILL_32_DFFSR_14 ( );
FILL FILL_33_DFFSR_14 ( );
FILL FILL_34_DFFSR_14 ( );
FILL FILL_35_DFFSR_14 ( );
FILL FILL_36_DFFSR_14 ( );
FILL FILL_37_DFFSR_14 ( );
FILL FILL_38_DFFSR_14 ( );
FILL FILL_39_DFFSR_14 ( );
FILL FILL_40_DFFSR_14 ( );
FILL FILL_41_DFFSR_14 ( );
FILL FILL_42_DFFSR_14 ( );
FILL FILL_43_DFFSR_14 ( );
FILL FILL_44_DFFSR_14 ( );
FILL FILL_45_DFFSR_14 ( );
FILL FILL_46_DFFSR_14 ( );
FILL FILL_47_DFFSR_14 ( );
FILL FILL_48_DFFSR_14 ( );
FILL FILL_49_DFFSR_14 ( );
FILL FILL_50_DFFSR_14 ( );
FILL FILL_51_DFFSR_14 ( );
FILL FILL_0_BUFX2_87 ( );
FILL FILL_1_BUFX2_87 ( );
FILL FILL_2_BUFX2_87 ( );
FILL FILL_3_BUFX2_87 ( );
FILL FILL_4_BUFX2_87 ( );
FILL FILL_5_BUFX2_87 ( );
FILL FILL_6_BUFX2_87 ( );
FILL FILL_0_CLKBUF1_26 ( );
FILL FILL_1_CLKBUF1_26 ( );
FILL FILL_2_CLKBUF1_26 ( );
FILL FILL_3_CLKBUF1_26 ( );
FILL FILL_4_CLKBUF1_26 ( );
FILL FILL_5_CLKBUF1_26 ( );
FILL FILL_6_CLKBUF1_26 ( );
FILL FILL_7_CLKBUF1_26 ( );
FILL FILL_8_CLKBUF1_26 ( );
FILL FILL_9_CLKBUF1_26 ( );
FILL FILL_10_CLKBUF1_26 ( );
FILL FILL_11_CLKBUF1_26 ( );
FILL FILL_12_CLKBUF1_26 ( );
FILL FILL_13_CLKBUF1_26 ( );
FILL FILL_14_CLKBUF1_26 ( );
FILL FILL_15_CLKBUF1_26 ( );
FILL FILL_16_CLKBUF1_26 ( );
FILL FILL_17_CLKBUF1_26 ( );
FILL FILL_18_CLKBUF1_26 ( );
FILL FILL_19_CLKBUF1_26 ( );
FILL FILL_20_CLKBUF1_26 ( );
FILL FILL_0_INVX1_31 ( );
FILL FILL_1_INVX1_31 ( );
FILL FILL_2_INVX1_31 ( );
FILL FILL_3_INVX1_31 ( );
FILL FILL_4_INVX1_31 ( );
FILL FILL_0_OAI22X1_13 ( );
FILL FILL_1_OAI22X1_13 ( );
FILL FILL_2_OAI22X1_13 ( );
FILL FILL_3_OAI22X1_13 ( );
FILL FILL_4_OAI22X1_13 ( );
FILL FILL_5_OAI22X1_13 ( );
FILL FILL_6_OAI22X1_13 ( );
FILL FILL_7_OAI22X1_13 ( );
FILL FILL_8_OAI22X1_13 ( );
FILL FILL_9_OAI22X1_13 ( );
FILL FILL_10_OAI22X1_13 ( );
FILL FILL_0_OAI22X1_1 ( );
FILL FILL_1_OAI22X1_1 ( );
FILL FILL_2_OAI22X1_1 ( );
FILL FILL_3_OAI22X1_1 ( );
FILL FILL_4_OAI22X1_1 ( );
FILL FILL_5_OAI22X1_1 ( );
FILL FILL_6_OAI22X1_1 ( );
FILL FILL_7_OAI22X1_1 ( );
FILL FILL_8_OAI22X1_1 ( );
FILL FILL_9_OAI22X1_1 ( );
FILL FILL_10_OAI22X1_1 ( );
FILL FILL_0_INVX1_1 ( );
FILL FILL_1_INVX1_1 ( );
FILL FILL_2_INVX1_1 ( );
FILL FILL_3_INVX1_1 ( );
FILL FILL_4_INVX1_1 ( );
FILL FILL_0_DFFSR_105 ( );
FILL FILL_1_DFFSR_105 ( );
FILL FILL_2_DFFSR_105 ( );
FILL FILL_3_DFFSR_105 ( );
FILL FILL_4_DFFSR_105 ( );
FILL FILL_5_DFFSR_105 ( );
FILL FILL_6_DFFSR_105 ( );
FILL FILL_7_DFFSR_105 ( );
FILL FILL_8_DFFSR_105 ( );
FILL FILL_9_DFFSR_105 ( );
FILL FILL_10_DFFSR_105 ( );
FILL FILL_11_DFFSR_105 ( );
FILL FILL_12_DFFSR_105 ( );
FILL FILL_13_DFFSR_105 ( );
FILL FILL_14_DFFSR_105 ( );
FILL FILL_15_DFFSR_105 ( );
FILL FILL_16_DFFSR_105 ( );
FILL FILL_17_DFFSR_105 ( );
FILL FILL_18_DFFSR_105 ( );
FILL FILL_19_DFFSR_105 ( );
FILL FILL_20_DFFSR_105 ( );
FILL FILL_21_DFFSR_105 ( );
FILL FILL_22_DFFSR_105 ( );
FILL FILL_23_DFFSR_105 ( );
FILL FILL_24_DFFSR_105 ( );
FILL FILL_25_DFFSR_105 ( );
FILL FILL_26_DFFSR_105 ( );
FILL FILL_27_DFFSR_105 ( );
FILL FILL_28_DFFSR_105 ( );
FILL FILL_29_DFFSR_105 ( );
FILL FILL_30_DFFSR_105 ( );
FILL FILL_31_DFFSR_105 ( );
FILL FILL_32_DFFSR_105 ( );
FILL FILL_33_DFFSR_105 ( );
FILL FILL_34_DFFSR_105 ( );
FILL FILL_35_DFFSR_105 ( );
FILL FILL_36_DFFSR_105 ( );
FILL FILL_37_DFFSR_105 ( );
FILL FILL_38_DFFSR_105 ( );
FILL FILL_39_DFFSR_105 ( );
FILL FILL_40_DFFSR_105 ( );
FILL FILL_41_DFFSR_105 ( );
FILL FILL_42_DFFSR_105 ( );
FILL FILL_43_DFFSR_105 ( );
FILL FILL_44_DFFSR_105 ( );
FILL FILL_45_DFFSR_105 ( );
FILL FILL_46_DFFSR_105 ( );
FILL FILL_47_DFFSR_105 ( );
FILL FILL_48_DFFSR_105 ( );
FILL FILL_49_DFFSR_105 ( );
FILL FILL_50_DFFSR_105 ( );
FILL FILL_51_DFFSR_105 ( );
FILL FILL_0_DFFSR_134 ( );
FILL FILL_1_DFFSR_134 ( );
FILL FILL_2_DFFSR_134 ( );
FILL FILL_3_DFFSR_134 ( );
FILL FILL_4_DFFSR_134 ( );
FILL FILL_5_DFFSR_134 ( );
FILL FILL_6_DFFSR_134 ( );
FILL FILL_7_DFFSR_134 ( );
FILL FILL_8_DFFSR_134 ( );
FILL FILL_9_DFFSR_134 ( );
FILL FILL_10_DFFSR_134 ( );
FILL FILL_11_DFFSR_134 ( );
FILL FILL_12_DFFSR_134 ( );
FILL FILL_13_DFFSR_134 ( );
FILL FILL_14_DFFSR_134 ( );
FILL FILL_15_DFFSR_134 ( );
FILL FILL_16_DFFSR_134 ( );
FILL FILL_17_DFFSR_134 ( );
FILL FILL_18_DFFSR_134 ( );
FILL FILL_19_DFFSR_134 ( );
FILL FILL_20_DFFSR_134 ( );
FILL FILL_21_DFFSR_134 ( );
FILL FILL_22_DFFSR_134 ( );
FILL FILL_23_DFFSR_134 ( );
FILL FILL_24_DFFSR_134 ( );
FILL FILL_25_DFFSR_134 ( );
FILL FILL_26_DFFSR_134 ( );
FILL FILL_27_DFFSR_134 ( );
FILL FILL_28_DFFSR_134 ( );
FILL FILL_29_DFFSR_134 ( );
FILL FILL_30_DFFSR_134 ( );
FILL FILL_31_DFFSR_134 ( );
FILL FILL_32_DFFSR_134 ( );
FILL FILL_33_DFFSR_134 ( );
FILL FILL_34_DFFSR_134 ( );
FILL FILL_35_DFFSR_134 ( );
FILL FILL_36_DFFSR_134 ( );
FILL FILL_37_DFFSR_134 ( );
FILL FILL_38_DFFSR_134 ( );
FILL FILL_39_DFFSR_134 ( );
FILL FILL_40_DFFSR_134 ( );
FILL FILL_41_DFFSR_134 ( );
FILL FILL_42_DFFSR_134 ( );
FILL FILL_43_DFFSR_134 ( );
FILL FILL_44_DFFSR_134 ( );
FILL FILL_45_DFFSR_134 ( );
FILL FILL_46_DFFSR_134 ( );
FILL FILL_47_DFFSR_134 ( );
FILL FILL_48_DFFSR_134 ( );
FILL FILL_49_DFFSR_134 ( );
FILL FILL_50_DFFSR_134 ( );
FILL FILL_51_DFFSR_134 ( );
FILL FILL_0_NAND3X1_76 ( );
FILL FILL_1_NAND3X1_76 ( );
FILL FILL_2_NAND3X1_76 ( );
FILL FILL_3_NAND3X1_76 ( );
FILL FILL_4_NAND3X1_76 ( );
FILL FILL_5_NAND3X1_76 ( );
FILL FILL_6_NAND3X1_76 ( );
FILL FILL_7_NAND3X1_76 ( );
FILL FILL_8_NAND3X1_76 ( );
FILL FILL_0_CLKBUF1_39 ( );
FILL FILL_1_CLKBUF1_39 ( );
FILL FILL_2_CLKBUF1_39 ( );
FILL FILL_3_CLKBUF1_39 ( );
FILL FILL_4_CLKBUF1_39 ( );
FILL FILL_5_CLKBUF1_39 ( );
FILL FILL_6_CLKBUF1_39 ( );
FILL FILL_7_CLKBUF1_39 ( );
FILL FILL_8_CLKBUF1_39 ( );
FILL FILL_9_CLKBUF1_39 ( );
FILL FILL_10_CLKBUF1_39 ( );
FILL FILL_11_CLKBUF1_39 ( );
FILL FILL_12_CLKBUF1_39 ( );
FILL FILL_13_CLKBUF1_39 ( );
FILL FILL_14_CLKBUF1_39 ( );
FILL FILL_15_CLKBUF1_39 ( );
FILL FILL_16_CLKBUF1_39 ( );
FILL FILL_17_CLKBUF1_39 ( );
FILL FILL_18_CLKBUF1_39 ( );
FILL FILL_19_CLKBUF1_39 ( );
FILL FILL_20_CLKBUF1_39 ( );
FILL FILL_0_DFFSR_152 ( );
FILL FILL_1_DFFSR_152 ( );
FILL FILL_2_DFFSR_152 ( );
FILL FILL_3_DFFSR_152 ( );
FILL FILL_4_DFFSR_152 ( );
FILL FILL_5_DFFSR_152 ( );
FILL FILL_6_DFFSR_152 ( );
FILL FILL_7_DFFSR_152 ( );
FILL FILL_8_DFFSR_152 ( );
FILL FILL_9_DFFSR_152 ( );
FILL FILL_10_DFFSR_152 ( );
FILL FILL_11_DFFSR_152 ( );
FILL FILL_12_DFFSR_152 ( );
FILL FILL_13_DFFSR_152 ( );
FILL FILL_14_DFFSR_152 ( );
FILL FILL_15_DFFSR_152 ( );
FILL FILL_16_DFFSR_152 ( );
FILL FILL_17_DFFSR_152 ( );
FILL FILL_18_DFFSR_152 ( );
FILL FILL_19_DFFSR_152 ( );
FILL FILL_20_DFFSR_152 ( );
FILL FILL_21_DFFSR_152 ( );
FILL FILL_22_DFFSR_152 ( );
FILL FILL_23_DFFSR_152 ( );
FILL FILL_24_DFFSR_152 ( );
FILL FILL_25_DFFSR_152 ( );
FILL FILL_26_DFFSR_152 ( );
FILL FILL_27_DFFSR_152 ( );
FILL FILL_28_DFFSR_152 ( );
FILL FILL_29_DFFSR_152 ( );
FILL FILL_30_DFFSR_152 ( );
FILL FILL_31_DFFSR_152 ( );
FILL FILL_32_DFFSR_152 ( );
FILL FILL_33_DFFSR_152 ( );
FILL FILL_34_DFFSR_152 ( );
FILL FILL_35_DFFSR_152 ( );
FILL FILL_36_DFFSR_152 ( );
FILL FILL_37_DFFSR_152 ( );
FILL FILL_38_DFFSR_152 ( );
FILL FILL_39_DFFSR_152 ( );
FILL FILL_40_DFFSR_152 ( );
FILL FILL_41_DFFSR_152 ( );
FILL FILL_42_DFFSR_152 ( );
FILL FILL_43_DFFSR_152 ( );
FILL FILL_44_DFFSR_152 ( );
FILL FILL_45_DFFSR_152 ( );
FILL FILL_46_DFFSR_152 ( );
FILL FILL_47_DFFSR_152 ( );
FILL FILL_48_DFFSR_152 ( );
FILL FILL_49_DFFSR_152 ( );
FILL FILL_50_DFFSR_152 ( );
FILL FILL_51_DFFSR_152 ( );
FILL FILL_0_NAND2X1_104 ( );
FILL FILL_1_NAND2X1_104 ( );
FILL FILL_2_NAND2X1_104 ( );
FILL FILL_3_NAND2X1_104 ( );
FILL FILL_4_NAND2X1_104 ( );
FILL FILL_5_NAND2X1_104 ( );
FILL FILL_6_NAND2X1_104 ( );
FILL FILL_0_NAND2X1_105 ( );
FILL FILL_1_NAND2X1_105 ( );
FILL FILL_2_NAND2X1_105 ( );
FILL FILL_3_NAND2X1_105 ( );
FILL FILL_4_NAND2X1_105 ( );
FILL FILL_5_NAND2X1_105 ( );
FILL FILL_6_NAND2X1_105 ( );
FILL FILL_0_NAND2X1_98 ( );
FILL FILL_1_NAND2X1_98 ( );
FILL FILL_2_NAND2X1_98 ( );
FILL FILL_3_NAND2X1_98 ( );
FILL FILL_4_NAND2X1_98 ( );
FILL FILL_5_NAND2X1_98 ( );
FILL FILL_6_NAND2X1_98 ( );
FILL FILL_0_AOI22X1_28 ( );
FILL FILL_1_AOI22X1_28 ( );
FILL FILL_2_AOI22X1_28 ( );
FILL FILL_3_AOI22X1_28 ( );
FILL FILL_4_AOI22X1_28 ( );
FILL FILL_5_AOI22X1_28 ( );
FILL FILL_6_AOI22X1_28 ( );
FILL FILL_7_AOI22X1_28 ( );
FILL FILL_8_AOI22X1_28 ( );
FILL FILL_9_AOI22X1_28 ( );
FILL FILL_10_AOI22X1_28 ( );
FILL FILL_11_AOI22X1_28 ( );
FILL FILL_0_NAND3X1_204 ( );
FILL FILL_1_NAND3X1_204 ( );
FILL FILL_2_NAND3X1_204 ( );
FILL FILL_3_NAND3X1_204 ( );
FILL FILL_4_NAND3X1_204 ( );
FILL FILL_5_NAND3X1_204 ( );
FILL FILL_6_NAND3X1_204 ( );
FILL FILL_7_NAND3X1_204 ( );
FILL FILL_8_NAND3X1_204 ( );
FILL FILL_9_NAND3X1_204 ( );
FILL FILL_0_NAND3X1_200 ( );
FILL FILL_1_NAND3X1_200 ( );
FILL FILL_2_NAND3X1_200 ( );
FILL FILL_3_NAND3X1_200 ( );
FILL FILL_4_NAND3X1_200 ( );
FILL FILL_5_NAND3X1_200 ( );
FILL FILL_6_NAND3X1_200 ( );
FILL FILL_7_NAND3X1_200 ( );
FILL FILL_8_NAND3X1_200 ( );
FILL FILL_0_INVX1_167 ( );
FILL FILL_1_INVX1_167 ( );
FILL FILL_2_INVX1_167 ( );
FILL FILL_3_INVX1_167 ( );
FILL FILL_4_INVX1_167 ( );
FILL FILL_0_NAND3X1_202 ( );
FILL FILL_1_NAND3X1_202 ( );
FILL FILL_2_NAND3X1_202 ( );
FILL FILL_3_NAND3X1_202 ( );
FILL FILL_4_NAND3X1_202 ( );
FILL FILL_5_NAND3X1_202 ( );
FILL FILL_6_NAND3X1_202 ( );
FILL FILL_7_NAND3X1_202 ( );
FILL FILL_8_NAND3X1_202 ( );
FILL FILL_9_NAND3X1_202 ( );
FILL FILL_0_NAND2X1_96 ( );
FILL FILL_1_NAND2X1_96 ( );
FILL FILL_2_NAND2X1_96 ( );
FILL FILL_3_NAND2X1_96 ( );
FILL FILL_4_NAND2X1_96 ( );
FILL FILL_5_NAND2X1_96 ( );
FILL FILL_6_NAND2X1_96 ( );
FILL FILL_0_NAND2X1_106 ( );
FILL FILL_1_NAND2X1_106 ( );
FILL FILL_2_NAND2X1_106 ( );
FILL FILL_3_NAND2X1_106 ( );
FILL FILL_4_NAND2X1_106 ( );
FILL FILL_5_NAND2X1_106 ( );
FILL FILL_6_NAND2X1_106 ( );
FILL FILL_0_AOI21X1_52 ( );
FILL FILL_1_AOI21X1_52 ( );
FILL FILL_2_AOI21X1_52 ( );
FILL FILL_3_AOI21X1_52 ( );
FILL FILL_4_AOI21X1_52 ( );
FILL FILL_5_AOI21X1_52 ( );
FILL FILL_6_AOI21X1_52 ( );
FILL FILL_7_AOI21X1_52 ( );
FILL FILL_8_AOI21X1_52 ( );
FILL FILL_0_DFFSR_280 ( );
FILL FILL_1_DFFSR_280 ( );
FILL FILL_2_DFFSR_280 ( );
FILL FILL_3_DFFSR_280 ( );
FILL FILL_4_DFFSR_280 ( );
FILL FILL_5_DFFSR_280 ( );
FILL FILL_6_DFFSR_280 ( );
FILL FILL_7_DFFSR_280 ( );
FILL FILL_8_DFFSR_280 ( );
FILL FILL_9_DFFSR_280 ( );
FILL FILL_10_DFFSR_280 ( );
FILL FILL_11_DFFSR_280 ( );
FILL FILL_12_DFFSR_280 ( );
FILL FILL_13_DFFSR_280 ( );
FILL FILL_14_DFFSR_280 ( );
FILL FILL_15_DFFSR_280 ( );
FILL FILL_16_DFFSR_280 ( );
FILL FILL_17_DFFSR_280 ( );
FILL FILL_18_DFFSR_280 ( );
FILL FILL_19_DFFSR_280 ( );
FILL FILL_20_DFFSR_280 ( );
FILL FILL_21_DFFSR_280 ( );
FILL FILL_22_DFFSR_280 ( );
FILL FILL_23_DFFSR_280 ( );
FILL FILL_24_DFFSR_280 ( );
FILL FILL_25_DFFSR_280 ( );
FILL FILL_26_DFFSR_280 ( );
FILL FILL_27_DFFSR_280 ( );
FILL FILL_28_DFFSR_280 ( );
FILL FILL_29_DFFSR_280 ( );
FILL FILL_30_DFFSR_280 ( );
FILL FILL_31_DFFSR_280 ( );
FILL FILL_32_DFFSR_280 ( );
FILL FILL_33_DFFSR_280 ( );
FILL FILL_34_DFFSR_280 ( );
FILL FILL_35_DFFSR_280 ( );
FILL FILL_36_DFFSR_280 ( );
FILL FILL_37_DFFSR_280 ( );
FILL FILL_38_DFFSR_280 ( );
FILL FILL_39_DFFSR_280 ( );
FILL FILL_40_DFFSR_280 ( );
FILL FILL_41_DFFSR_280 ( );
FILL FILL_42_DFFSR_280 ( );
FILL FILL_43_DFFSR_280 ( );
FILL FILL_44_DFFSR_280 ( );
FILL FILL_45_DFFSR_280 ( );
FILL FILL_46_DFFSR_280 ( );
FILL FILL_47_DFFSR_280 ( );
FILL FILL_48_DFFSR_280 ( );
FILL FILL_49_DFFSR_280 ( );
FILL FILL_50_DFFSR_280 ( );
FILL FILL_0_NOR2X1_5 ( );
FILL FILL_1_NOR2X1_5 ( );
FILL FILL_2_NOR2X1_5 ( );
FILL FILL_3_NOR2X1_5 ( );
FILL FILL_4_NOR2X1_5 ( );
FILL FILL_5_NOR2X1_5 ( );
FILL FILL_6_NOR2X1_5 ( );
FILL FILL_0_NAND2X1_7 ( );
FILL FILL_1_NAND2X1_7 ( );
FILL FILL_2_NAND2X1_7 ( );
FILL FILL_3_NAND2X1_7 ( );
FILL FILL_4_NAND2X1_7 ( );
FILL FILL_5_NAND2X1_7 ( );
FILL FILL_6_NAND2X1_7 ( );
FILL FILL_0_OAI21X1_118 ( );
FILL FILL_1_OAI21X1_118 ( );
FILL FILL_2_OAI21X1_118 ( );
FILL FILL_3_OAI21X1_118 ( );
FILL FILL_4_OAI21X1_118 ( );
FILL FILL_5_OAI21X1_118 ( );
FILL FILL_6_OAI21X1_118 ( );
FILL FILL_7_OAI21X1_118 ( );
FILL FILL_8_OAI21X1_118 ( );
FILL FILL_0_OR2X2_6 ( );
FILL FILL_1_OR2X2_6 ( );
FILL FILL_2_OR2X2_6 ( );
FILL FILL_3_OR2X2_6 ( );
FILL FILL_4_OR2X2_6 ( );
FILL FILL_5_OR2X2_6 ( );
FILL FILL_6_OR2X2_6 ( );
FILL FILL_7_OR2X2_6 ( );
FILL FILL_8_OR2X2_6 ( );
FILL FILL_9_OR2X2_6 ( );
FILL FILL_0_OAI21X1_119 ( );
FILL FILL_1_OAI21X1_119 ( );
FILL FILL_2_OAI21X1_119 ( );
FILL FILL_3_OAI21X1_119 ( );
FILL FILL_4_OAI21X1_119 ( );
FILL FILL_5_OAI21X1_119 ( );
FILL FILL_6_OAI21X1_119 ( );
FILL FILL_7_OAI21X1_119 ( );
FILL FILL_8_OAI21X1_119 ( );
FILL FILL_0_OAI21X1_4 ( );
FILL FILL_1_OAI21X1_4 ( );
FILL FILL_2_OAI21X1_4 ( );
FILL FILL_3_OAI21X1_4 ( );
FILL FILL_4_OAI21X1_4 ( );
FILL FILL_5_OAI21X1_4 ( );
FILL FILL_6_OAI21X1_4 ( );
FILL FILL_7_OAI21X1_4 ( );
FILL FILL_8_OAI21X1_4 ( );
FILL FILL_9_OAI21X1_4 ( );
FILL FILL_0_NAND3X1_22 ( );
FILL FILL_1_NAND3X1_22 ( );
FILL FILL_2_NAND3X1_22 ( );
FILL FILL_3_NAND3X1_22 ( );
FILL FILL_4_NAND3X1_22 ( );
FILL FILL_5_NAND3X1_22 ( );
FILL FILL_6_NAND3X1_22 ( );
FILL FILL_7_NAND3X1_22 ( );
FILL FILL_8_NAND3X1_22 ( );
FILL FILL_0_INVX1_49 ( );
FILL FILL_1_INVX1_49 ( );
FILL FILL_2_INVX1_49 ( );
FILL FILL_3_INVX1_49 ( );
FILL FILL_0_NAND3X1_23 ( );
FILL FILL_1_NAND3X1_23 ( );
FILL FILL_2_NAND3X1_23 ( );
FILL FILL_3_NAND3X1_23 ( );
FILL FILL_4_NAND3X1_23 ( );
FILL FILL_5_NAND3X1_23 ( );
FILL FILL_6_NAND3X1_23 ( );
FILL FILL_7_NAND3X1_23 ( );
FILL FILL_8_NAND3X1_23 ( );
FILL FILL_0_NAND3X1_21 ( );
FILL FILL_1_NAND3X1_21 ( );
FILL FILL_2_NAND3X1_21 ( );
FILL FILL_3_NAND3X1_21 ( );
FILL FILL_4_NAND3X1_21 ( );
FILL FILL_5_NAND3X1_21 ( );
FILL FILL_6_NAND3X1_21 ( );
FILL FILL_7_NAND3X1_21 ( );
FILL FILL_8_NAND3X1_21 ( );
FILL FILL_0_BUFX2_22 ( );
FILL FILL_1_BUFX2_22 ( );
FILL FILL_2_BUFX2_22 ( );
FILL FILL_3_BUFX2_22 ( );
FILL FILL_4_BUFX2_22 ( );
FILL FILL_5_BUFX2_22 ( );
FILL FILL_6_BUFX2_22 ( );
FILL FILL_0_DFFSR_13 ( );
FILL FILL_1_DFFSR_13 ( );
FILL FILL_2_DFFSR_13 ( );
FILL FILL_3_DFFSR_13 ( );
FILL FILL_4_DFFSR_13 ( );
FILL FILL_5_DFFSR_13 ( );
FILL FILL_6_DFFSR_13 ( );
FILL FILL_7_DFFSR_13 ( );
FILL FILL_8_DFFSR_13 ( );
FILL FILL_9_DFFSR_13 ( );
FILL FILL_10_DFFSR_13 ( );
FILL FILL_11_DFFSR_13 ( );
FILL FILL_12_DFFSR_13 ( );
FILL FILL_13_DFFSR_13 ( );
FILL FILL_14_DFFSR_13 ( );
FILL FILL_15_DFFSR_13 ( );
FILL FILL_16_DFFSR_13 ( );
FILL FILL_17_DFFSR_13 ( );
FILL FILL_18_DFFSR_13 ( );
FILL FILL_19_DFFSR_13 ( );
FILL FILL_20_DFFSR_13 ( );
FILL FILL_21_DFFSR_13 ( );
FILL FILL_22_DFFSR_13 ( );
FILL FILL_23_DFFSR_13 ( );
FILL FILL_24_DFFSR_13 ( );
FILL FILL_25_DFFSR_13 ( );
FILL FILL_26_DFFSR_13 ( );
FILL FILL_27_DFFSR_13 ( );
FILL FILL_28_DFFSR_13 ( );
FILL FILL_29_DFFSR_13 ( );
FILL FILL_30_DFFSR_13 ( );
FILL FILL_31_DFFSR_13 ( );
FILL FILL_32_DFFSR_13 ( );
FILL FILL_33_DFFSR_13 ( );
FILL FILL_34_DFFSR_13 ( );
FILL FILL_35_DFFSR_13 ( );
FILL FILL_36_DFFSR_13 ( );
FILL FILL_37_DFFSR_13 ( );
FILL FILL_38_DFFSR_13 ( );
FILL FILL_39_DFFSR_13 ( );
FILL FILL_40_DFFSR_13 ( );
FILL FILL_41_DFFSR_13 ( );
FILL FILL_42_DFFSR_13 ( );
FILL FILL_43_DFFSR_13 ( );
FILL FILL_44_DFFSR_13 ( );
FILL FILL_45_DFFSR_13 ( );
FILL FILL_46_DFFSR_13 ( );
FILL FILL_47_DFFSR_13 ( );
FILL FILL_48_DFFSR_13 ( );
FILL FILL_49_DFFSR_13 ( );
FILL FILL_50_DFFSR_13 ( );
FILL FILL_0_INVX1_32 ( );
FILL FILL_1_INVX1_32 ( );
FILL FILL_2_INVX1_32 ( );
FILL FILL_3_INVX1_32 ( );
FILL FILL_4_INVX1_32 ( );
FILL FILL_0_DFFSR_53 ( );
FILL FILL_1_DFFSR_53 ( );
FILL FILL_2_DFFSR_53 ( );
FILL FILL_3_DFFSR_53 ( );
FILL FILL_4_DFFSR_53 ( );
FILL FILL_5_DFFSR_53 ( );
FILL FILL_6_DFFSR_53 ( );
FILL FILL_7_DFFSR_53 ( );
FILL FILL_8_DFFSR_53 ( );
FILL FILL_9_DFFSR_53 ( );
FILL FILL_10_DFFSR_53 ( );
FILL FILL_11_DFFSR_53 ( );
FILL FILL_12_DFFSR_53 ( );
FILL FILL_13_DFFSR_53 ( );
FILL FILL_14_DFFSR_53 ( );
FILL FILL_15_DFFSR_53 ( );
FILL FILL_16_DFFSR_53 ( );
FILL FILL_17_DFFSR_53 ( );
FILL FILL_18_DFFSR_53 ( );
FILL FILL_19_DFFSR_53 ( );
FILL FILL_20_DFFSR_53 ( );
FILL FILL_21_DFFSR_53 ( );
FILL FILL_22_DFFSR_53 ( );
FILL FILL_23_DFFSR_53 ( );
FILL FILL_24_DFFSR_53 ( );
FILL FILL_25_DFFSR_53 ( );
FILL FILL_26_DFFSR_53 ( );
FILL FILL_27_DFFSR_53 ( );
FILL FILL_28_DFFSR_53 ( );
FILL FILL_29_DFFSR_53 ( );
FILL FILL_30_DFFSR_53 ( );
FILL FILL_31_DFFSR_53 ( );
FILL FILL_32_DFFSR_53 ( );
FILL FILL_33_DFFSR_53 ( );
FILL FILL_34_DFFSR_53 ( );
FILL FILL_35_DFFSR_53 ( );
FILL FILL_36_DFFSR_53 ( );
FILL FILL_37_DFFSR_53 ( );
FILL FILL_38_DFFSR_53 ( );
FILL FILL_39_DFFSR_53 ( );
FILL FILL_40_DFFSR_53 ( );
FILL FILL_41_DFFSR_53 ( );
FILL FILL_42_DFFSR_53 ( );
FILL FILL_43_DFFSR_53 ( );
FILL FILL_44_DFFSR_53 ( );
FILL FILL_45_DFFSR_53 ( );
FILL FILL_46_DFFSR_53 ( );
FILL FILL_47_DFFSR_53 ( );
FILL FILL_48_DFFSR_53 ( );
FILL FILL_49_DFFSR_53 ( );
FILL FILL_50_DFFSR_53 ( );
FILL FILL_0_DFFSR_121 ( );
FILL FILL_1_DFFSR_121 ( );
FILL FILL_2_DFFSR_121 ( );
FILL FILL_3_DFFSR_121 ( );
FILL FILL_4_DFFSR_121 ( );
FILL FILL_5_DFFSR_121 ( );
FILL FILL_6_DFFSR_121 ( );
FILL FILL_7_DFFSR_121 ( );
FILL FILL_8_DFFSR_121 ( );
FILL FILL_9_DFFSR_121 ( );
FILL FILL_10_DFFSR_121 ( );
FILL FILL_11_DFFSR_121 ( );
FILL FILL_12_DFFSR_121 ( );
FILL FILL_13_DFFSR_121 ( );
FILL FILL_14_DFFSR_121 ( );
FILL FILL_15_DFFSR_121 ( );
FILL FILL_16_DFFSR_121 ( );
FILL FILL_17_DFFSR_121 ( );
FILL FILL_18_DFFSR_121 ( );
FILL FILL_19_DFFSR_121 ( );
FILL FILL_20_DFFSR_121 ( );
FILL FILL_21_DFFSR_121 ( );
FILL FILL_22_DFFSR_121 ( );
FILL FILL_23_DFFSR_121 ( );
FILL FILL_24_DFFSR_121 ( );
FILL FILL_25_DFFSR_121 ( );
FILL FILL_26_DFFSR_121 ( );
FILL FILL_27_DFFSR_121 ( );
FILL FILL_28_DFFSR_121 ( );
FILL FILL_29_DFFSR_121 ( );
FILL FILL_30_DFFSR_121 ( );
FILL FILL_31_DFFSR_121 ( );
FILL FILL_32_DFFSR_121 ( );
FILL FILL_33_DFFSR_121 ( );
FILL FILL_34_DFFSR_121 ( );
FILL FILL_35_DFFSR_121 ( );
FILL FILL_36_DFFSR_121 ( );
FILL FILL_37_DFFSR_121 ( );
FILL FILL_38_DFFSR_121 ( );
FILL FILL_39_DFFSR_121 ( );
FILL FILL_40_DFFSR_121 ( );
FILL FILL_41_DFFSR_121 ( );
FILL FILL_42_DFFSR_121 ( );
FILL FILL_43_DFFSR_121 ( );
FILL FILL_44_DFFSR_121 ( );
FILL FILL_45_DFFSR_121 ( );
FILL FILL_46_DFFSR_121 ( );
FILL FILL_47_DFFSR_121 ( );
FILL FILL_48_DFFSR_121 ( );
FILL FILL_49_DFFSR_121 ( );
FILL FILL_50_DFFSR_121 ( );
FILL FILL_0_NAND2X1_40 ( );
FILL FILL_1_NAND2X1_40 ( );
FILL FILL_2_NAND2X1_40 ( );
FILL FILL_3_NAND2X1_40 ( );
FILL FILL_4_NAND2X1_40 ( );
FILL FILL_5_NAND2X1_40 ( );
FILL FILL_6_NAND2X1_40 ( );
FILL FILL_0_AND2X2_20 ( );
FILL FILL_1_AND2X2_20 ( );
FILL FILL_2_AND2X2_20 ( );
FILL FILL_3_AND2X2_20 ( );
FILL FILL_4_AND2X2_20 ( );
FILL FILL_5_AND2X2_20 ( );
FILL FILL_6_AND2X2_20 ( );
FILL FILL_7_AND2X2_20 ( );
FILL FILL_8_AND2X2_20 ( );
FILL FILL_9_AND2X2_20 ( );
FILL FILL_0_INVX1_110 ( );
FILL FILL_1_INVX1_110 ( );
FILL FILL_2_INVX1_110 ( );
FILL FILL_3_INVX1_110 ( );
FILL FILL_0_NAND2X1_52 ( );
FILL FILL_1_NAND2X1_52 ( );
FILL FILL_2_NAND2X1_52 ( );
FILL FILL_3_NAND2X1_52 ( );
FILL FILL_4_NAND2X1_52 ( );
FILL FILL_5_NAND2X1_52 ( );
FILL FILL_6_NAND2X1_52 ( );
FILL FILL_0_OAI22X1_30 ( );
FILL FILL_1_OAI22X1_30 ( );
FILL FILL_2_OAI22X1_30 ( );
FILL FILL_3_OAI22X1_30 ( );
FILL FILL_4_OAI22X1_30 ( );
FILL FILL_5_OAI22X1_30 ( );
FILL FILL_6_OAI22X1_30 ( );
FILL FILL_7_OAI22X1_30 ( );
FILL FILL_8_OAI22X1_30 ( );
FILL FILL_9_OAI22X1_30 ( );
FILL FILL_10_OAI22X1_30 ( );
FILL FILL_0_DFFSR_176 ( );
FILL FILL_1_DFFSR_176 ( );
FILL FILL_2_DFFSR_176 ( );
FILL FILL_3_DFFSR_176 ( );
FILL FILL_4_DFFSR_176 ( );
FILL FILL_5_DFFSR_176 ( );
FILL FILL_6_DFFSR_176 ( );
FILL FILL_7_DFFSR_176 ( );
FILL FILL_8_DFFSR_176 ( );
FILL FILL_9_DFFSR_176 ( );
FILL FILL_10_DFFSR_176 ( );
FILL FILL_11_DFFSR_176 ( );
FILL FILL_12_DFFSR_176 ( );
FILL FILL_13_DFFSR_176 ( );
FILL FILL_14_DFFSR_176 ( );
FILL FILL_15_DFFSR_176 ( );
FILL FILL_16_DFFSR_176 ( );
FILL FILL_17_DFFSR_176 ( );
FILL FILL_18_DFFSR_176 ( );
FILL FILL_19_DFFSR_176 ( );
FILL FILL_20_DFFSR_176 ( );
FILL FILL_21_DFFSR_176 ( );
FILL FILL_22_DFFSR_176 ( );
FILL FILL_23_DFFSR_176 ( );
FILL FILL_24_DFFSR_176 ( );
FILL FILL_25_DFFSR_176 ( );
FILL FILL_26_DFFSR_176 ( );
FILL FILL_27_DFFSR_176 ( );
FILL FILL_28_DFFSR_176 ( );
FILL FILL_29_DFFSR_176 ( );
FILL FILL_30_DFFSR_176 ( );
FILL FILL_31_DFFSR_176 ( );
FILL FILL_32_DFFSR_176 ( );
FILL FILL_33_DFFSR_176 ( );
FILL FILL_34_DFFSR_176 ( );
FILL FILL_35_DFFSR_176 ( );
FILL FILL_36_DFFSR_176 ( );
FILL FILL_37_DFFSR_176 ( );
FILL FILL_38_DFFSR_176 ( );
FILL FILL_39_DFFSR_176 ( );
FILL FILL_40_DFFSR_176 ( );
FILL FILL_41_DFFSR_176 ( );
FILL FILL_42_DFFSR_176 ( );
FILL FILL_43_DFFSR_176 ( );
FILL FILL_44_DFFSR_176 ( );
FILL FILL_45_DFFSR_176 ( );
FILL FILL_46_DFFSR_176 ( );
FILL FILL_47_DFFSR_176 ( );
FILL FILL_48_DFFSR_176 ( );
FILL FILL_49_DFFSR_176 ( );
FILL FILL_50_DFFSR_176 ( );
FILL FILL_51_DFFSR_176 ( );
FILL FILL_0_XOR2X1_5 ( );
FILL FILL_1_XOR2X1_5 ( );
FILL FILL_2_XOR2X1_5 ( );
FILL FILL_3_XOR2X1_5 ( );
FILL FILL_4_XOR2X1_5 ( );
FILL FILL_5_XOR2X1_5 ( );
FILL FILL_6_XOR2X1_5 ( );
FILL FILL_7_XOR2X1_5 ( );
FILL FILL_8_XOR2X1_5 ( );
FILL FILL_9_XOR2X1_5 ( );
FILL FILL_10_XOR2X1_5 ( );
FILL FILL_11_XOR2X1_5 ( );
FILL FILL_12_XOR2X1_5 ( );
FILL FILL_13_XOR2X1_5 ( );
FILL FILL_14_XOR2X1_5 ( );
FILL FILL_15_XOR2X1_5 ( );
FILL FILL_0_NAND2X1_94 ( );
FILL FILL_1_NAND2X1_94 ( );
FILL FILL_2_NAND2X1_94 ( );
FILL FILL_3_NAND2X1_94 ( );
FILL FILL_4_NAND2X1_94 ( );
FILL FILL_5_NAND2X1_94 ( );
FILL FILL_6_NAND2X1_94 ( );
FILL FILL_0_NOR2X1_69 ( );
FILL FILL_1_NOR2X1_69 ( );
FILL FILL_2_NOR2X1_69 ( );
FILL FILL_3_NOR2X1_69 ( );
FILL FILL_4_NOR2X1_69 ( );
FILL FILL_5_NOR2X1_69 ( );
FILL FILL_6_NOR2X1_69 ( );
FILL FILL_0_OAI21X1_68 ( );
FILL FILL_1_OAI21X1_68 ( );
FILL FILL_2_OAI21X1_68 ( );
FILL FILL_3_OAI21X1_68 ( );
FILL FILL_4_OAI21X1_68 ( );
FILL FILL_5_OAI21X1_68 ( );
FILL FILL_6_OAI21X1_68 ( );
FILL FILL_7_OAI21X1_68 ( );
FILL FILL_8_OAI21X1_68 ( );
FILL FILL_0_AOI22X1_27 ( );
FILL FILL_1_AOI22X1_27 ( );
FILL FILL_2_AOI22X1_27 ( );
FILL FILL_3_AOI22X1_27 ( );
FILL FILL_4_AOI22X1_27 ( );
FILL FILL_5_AOI22X1_27 ( );
FILL FILL_6_AOI22X1_27 ( );
FILL FILL_7_AOI22X1_27 ( );
FILL FILL_8_AOI22X1_27 ( );
FILL FILL_9_AOI22X1_27 ( );
FILL FILL_10_AOI22X1_27 ( );
FILL FILL_11_AOI22X1_27 ( );
FILL FILL_0_BUFX2_73 ( );
FILL FILL_1_BUFX2_73 ( );
FILL FILL_2_BUFX2_73 ( );
FILL FILL_3_BUFX2_73 ( );
FILL FILL_4_BUFX2_73 ( );
FILL FILL_5_BUFX2_73 ( );
FILL FILL_6_BUFX2_73 ( );
FILL FILL_0_INVX1_168 ( );
FILL FILL_1_INVX1_168 ( );
FILL FILL_2_INVX1_168 ( );
FILL FILL_3_INVX1_168 ( );
FILL FILL_4_INVX1_168 ( );
FILL FILL_0_OAI21X1_78 ( );
FILL FILL_1_OAI21X1_78 ( );
FILL FILL_2_OAI21X1_78 ( );
FILL FILL_3_OAI21X1_78 ( );
FILL FILL_4_OAI21X1_78 ( );
FILL FILL_5_OAI21X1_78 ( );
FILL FILL_6_OAI21X1_78 ( );
FILL FILL_7_OAI21X1_78 ( );
FILL FILL_8_OAI21X1_78 ( );
FILL FILL_9_OAI21X1_78 ( );
FILL FILL_0_INVX1_201 ( );
FILL FILL_1_INVX1_201 ( );
FILL FILL_2_INVX1_201 ( );
FILL FILL_3_INVX1_201 ( );
FILL FILL_4_INVX1_201 ( );
FILL FILL_0_OAI21X1_103 ( );
FILL FILL_1_OAI21X1_103 ( );
FILL FILL_2_OAI21X1_103 ( );
FILL FILL_3_OAI21X1_103 ( );
FILL FILL_4_OAI21X1_103 ( );
FILL FILL_5_OAI21X1_103 ( );
FILL FILL_6_OAI21X1_103 ( );
FILL FILL_7_OAI21X1_103 ( );
FILL FILL_8_OAI21X1_103 ( );
FILL FILL_0_OAI21X1_107 ( );
FILL FILL_1_OAI21X1_107 ( );
FILL FILL_2_OAI21X1_107 ( );
FILL FILL_3_OAI21X1_107 ( );
FILL FILL_4_OAI21X1_107 ( );
FILL FILL_5_OAI21X1_107 ( );
FILL FILL_6_OAI21X1_107 ( );
FILL FILL_7_OAI21X1_107 ( );
FILL FILL_8_OAI21X1_107 ( );
FILL FILL_0_NAND2X1_138 ( );
FILL FILL_1_NAND2X1_138 ( );
FILL FILL_2_NAND2X1_138 ( );
FILL FILL_3_NAND2X1_138 ( );
FILL FILL_4_NAND2X1_138 ( );
FILL FILL_5_NAND2X1_138 ( );
FILL FILL_6_NAND2X1_138 ( );
FILL FILL_0_DFFSR_108 ( );
FILL FILL_1_DFFSR_108 ( );
FILL FILL_2_DFFSR_108 ( );
FILL FILL_3_DFFSR_108 ( );
FILL FILL_4_DFFSR_108 ( );
FILL FILL_5_DFFSR_108 ( );
FILL FILL_6_DFFSR_108 ( );
FILL FILL_7_DFFSR_108 ( );
FILL FILL_8_DFFSR_108 ( );
FILL FILL_9_DFFSR_108 ( );
FILL FILL_10_DFFSR_108 ( );
FILL FILL_11_DFFSR_108 ( );
FILL FILL_12_DFFSR_108 ( );
FILL FILL_13_DFFSR_108 ( );
FILL FILL_14_DFFSR_108 ( );
FILL FILL_15_DFFSR_108 ( );
FILL FILL_16_DFFSR_108 ( );
FILL FILL_17_DFFSR_108 ( );
FILL FILL_18_DFFSR_108 ( );
FILL FILL_19_DFFSR_108 ( );
FILL FILL_20_DFFSR_108 ( );
FILL FILL_21_DFFSR_108 ( );
FILL FILL_22_DFFSR_108 ( );
FILL FILL_23_DFFSR_108 ( );
FILL FILL_24_DFFSR_108 ( );
FILL FILL_25_DFFSR_108 ( );
FILL FILL_26_DFFSR_108 ( );
FILL FILL_27_DFFSR_108 ( );
FILL FILL_28_DFFSR_108 ( );
FILL FILL_29_DFFSR_108 ( );
FILL FILL_30_DFFSR_108 ( );
FILL FILL_31_DFFSR_108 ( );
FILL FILL_32_DFFSR_108 ( );
FILL FILL_33_DFFSR_108 ( );
FILL FILL_34_DFFSR_108 ( );
FILL FILL_35_DFFSR_108 ( );
FILL FILL_36_DFFSR_108 ( );
FILL FILL_37_DFFSR_108 ( );
FILL FILL_38_DFFSR_108 ( );
FILL FILL_39_DFFSR_108 ( );
FILL FILL_40_DFFSR_108 ( );
FILL FILL_41_DFFSR_108 ( );
FILL FILL_42_DFFSR_108 ( );
FILL FILL_43_DFFSR_108 ( );
FILL FILL_44_DFFSR_108 ( );
FILL FILL_45_DFFSR_108 ( );
FILL FILL_46_DFFSR_108 ( );
FILL FILL_47_DFFSR_108 ( );
FILL FILL_48_DFFSR_108 ( );
FILL FILL_49_DFFSR_108 ( );
FILL FILL_50_DFFSR_108 ( );
FILL FILL_51_DFFSR_108 ( );
FILL FILL_0_INVX1_26 ( );
FILL FILL_1_INVX1_26 ( );
FILL FILL_2_INVX1_26 ( );
FILL FILL_3_INVX1_26 ( );
FILL FILL_0_AOI21X1_70 ( );
FILL FILL_1_AOI21X1_70 ( );
FILL FILL_2_AOI21X1_70 ( );
FILL FILL_3_AOI21X1_70 ( );
FILL FILL_4_AOI21X1_70 ( );
FILL FILL_5_AOI21X1_70 ( );
FILL FILL_6_AOI21X1_70 ( );
FILL FILL_7_AOI21X1_70 ( );
FILL FILL_8_AOI21X1_70 ( );
FILL FILL_9_AOI21X1_70 ( );
FILL FILL_0_NOR2X1_83 ( );
FILL FILL_1_NOR2X1_83 ( );
FILL FILL_2_NOR2X1_83 ( );
FILL FILL_3_NOR2X1_83 ( );
FILL FILL_4_NOR2X1_83 ( );
FILL FILL_5_NOR2X1_83 ( );
FILL FILL_6_NOR2X1_83 ( );
FILL FILL_0_NAND2X1_182 ( );
FILL FILL_1_NAND2X1_182 ( );
FILL FILL_2_NAND2X1_182 ( );
FILL FILL_3_NAND2X1_182 ( );
FILL FILL_4_NAND2X1_182 ( );
FILL FILL_5_NAND2X1_182 ( );
FILL FILL_6_NAND2X1_182 ( );
FILL FILL_0_NAND3X1_249 ( );
FILL FILL_1_NAND3X1_249 ( );
FILL FILL_2_NAND3X1_249 ( );
FILL FILL_3_NAND3X1_249 ( );
FILL FILL_4_NAND3X1_249 ( );
FILL FILL_5_NAND3X1_249 ( );
FILL FILL_6_NAND3X1_249 ( );
FILL FILL_7_NAND3X1_249 ( );
FILL FILL_8_NAND3X1_249 ( );
FILL FILL_0_NAND2X1_17 ( );
FILL FILL_1_NAND2X1_17 ( );
FILL FILL_2_NAND2X1_17 ( );
FILL FILL_3_NAND2X1_17 ( );
FILL FILL_4_NAND2X1_17 ( );
FILL FILL_5_NAND2X1_17 ( );
FILL FILL_6_NAND2X1_17 ( );
FILL FILL_0_NAND3X1_41 ( );
FILL FILL_1_NAND3X1_41 ( );
FILL FILL_2_NAND3X1_41 ( );
FILL FILL_3_NAND3X1_41 ( );
FILL FILL_4_NAND3X1_41 ( );
FILL FILL_5_NAND3X1_41 ( );
FILL FILL_6_NAND3X1_41 ( );
FILL FILL_7_NAND3X1_41 ( );
FILL FILL_8_NAND3X1_41 ( );
FILL FILL_0_BUFX2_11 ( );
FILL FILL_1_BUFX2_11 ( );
FILL FILL_2_BUFX2_11 ( );
FILL FILL_3_BUFX2_11 ( );
FILL FILL_4_BUFX2_11 ( );
FILL FILL_5_BUFX2_11 ( );
FILL FILL_6_BUFX2_11 ( );
FILL FILL_7_BUFX2_11 ( );
FILL FILL_0_BUFX2_4 ( );
FILL FILL_1_BUFX2_4 ( );
FILL FILL_2_BUFX2_4 ( );
FILL FILL_3_BUFX2_4 ( );
FILL FILL_4_BUFX2_4 ( );
FILL FILL_5_BUFX2_4 ( );
FILL FILL_6_BUFX2_4 ( );
FILL FILL_0_DFFSR_107 ( );
FILL FILL_1_DFFSR_107 ( );
FILL FILL_2_DFFSR_107 ( );
FILL FILL_3_DFFSR_107 ( );
FILL FILL_4_DFFSR_107 ( );
FILL FILL_5_DFFSR_107 ( );
FILL FILL_6_DFFSR_107 ( );
FILL FILL_7_DFFSR_107 ( );
FILL FILL_8_DFFSR_107 ( );
FILL FILL_9_DFFSR_107 ( );
FILL FILL_10_DFFSR_107 ( );
FILL FILL_11_DFFSR_107 ( );
FILL FILL_12_DFFSR_107 ( );
FILL FILL_13_DFFSR_107 ( );
FILL FILL_14_DFFSR_107 ( );
FILL FILL_15_DFFSR_107 ( );
FILL FILL_16_DFFSR_107 ( );
FILL FILL_17_DFFSR_107 ( );
FILL FILL_18_DFFSR_107 ( );
FILL FILL_19_DFFSR_107 ( );
FILL FILL_20_DFFSR_107 ( );
FILL FILL_21_DFFSR_107 ( );
FILL FILL_22_DFFSR_107 ( );
FILL FILL_23_DFFSR_107 ( );
FILL FILL_24_DFFSR_107 ( );
FILL FILL_25_DFFSR_107 ( );
FILL FILL_26_DFFSR_107 ( );
FILL FILL_27_DFFSR_107 ( );
FILL FILL_28_DFFSR_107 ( );
FILL FILL_29_DFFSR_107 ( );
FILL FILL_30_DFFSR_107 ( );
FILL FILL_31_DFFSR_107 ( );
FILL FILL_32_DFFSR_107 ( );
FILL FILL_33_DFFSR_107 ( );
FILL FILL_34_DFFSR_107 ( );
FILL FILL_35_DFFSR_107 ( );
FILL FILL_36_DFFSR_107 ( );
FILL FILL_37_DFFSR_107 ( );
FILL FILL_38_DFFSR_107 ( );
FILL FILL_39_DFFSR_107 ( );
FILL FILL_40_DFFSR_107 ( );
FILL FILL_41_DFFSR_107 ( );
FILL FILL_42_DFFSR_107 ( );
FILL FILL_43_DFFSR_107 ( );
FILL FILL_44_DFFSR_107 ( );
FILL FILL_45_DFFSR_107 ( );
FILL FILL_46_DFFSR_107 ( );
FILL FILL_47_DFFSR_107 ( );
FILL FILL_48_DFFSR_107 ( );
FILL FILL_49_DFFSR_107 ( );
FILL FILL_50_DFFSR_107 ( );
FILL FILL_0_NAND3X1_7 ( );
FILL FILL_1_NAND3X1_7 ( );
FILL FILL_2_NAND3X1_7 ( );
FILL FILL_3_NAND3X1_7 ( );
FILL FILL_4_NAND3X1_7 ( );
FILL FILL_5_NAND3X1_7 ( );
FILL FILL_6_NAND3X1_7 ( );
FILL FILL_7_NAND3X1_7 ( );
FILL FILL_8_NAND3X1_7 ( );
FILL FILL_0_NOR2X1_8 ( );
FILL FILL_1_NOR2X1_8 ( );
FILL FILL_2_NOR2X1_8 ( );
FILL FILL_3_NOR2X1_8 ( );
FILL FILL_4_NOR2X1_8 ( );
FILL FILL_5_NOR2X1_8 ( );
FILL FILL_6_NOR2X1_8 ( );
FILL FILL_0_INVX1_2 ( );
FILL FILL_1_INVX1_2 ( );
FILL FILL_2_INVX1_2 ( );
FILL FILL_3_INVX1_2 ( );
FILL FILL_4_INVX1_2 ( );
FILL FILL_0_DFFSR_49 ( );
FILL FILL_1_DFFSR_49 ( );
FILL FILL_2_DFFSR_49 ( );
FILL FILL_3_DFFSR_49 ( );
FILL FILL_4_DFFSR_49 ( );
FILL FILL_5_DFFSR_49 ( );
FILL FILL_6_DFFSR_49 ( );
FILL FILL_7_DFFSR_49 ( );
FILL FILL_8_DFFSR_49 ( );
FILL FILL_9_DFFSR_49 ( );
FILL FILL_10_DFFSR_49 ( );
FILL FILL_11_DFFSR_49 ( );
FILL FILL_12_DFFSR_49 ( );
FILL FILL_13_DFFSR_49 ( );
FILL FILL_14_DFFSR_49 ( );
FILL FILL_15_DFFSR_49 ( );
FILL FILL_16_DFFSR_49 ( );
FILL FILL_17_DFFSR_49 ( );
FILL FILL_18_DFFSR_49 ( );
FILL FILL_19_DFFSR_49 ( );
FILL FILL_20_DFFSR_49 ( );
FILL FILL_21_DFFSR_49 ( );
FILL FILL_22_DFFSR_49 ( );
FILL FILL_23_DFFSR_49 ( );
FILL FILL_24_DFFSR_49 ( );
FILL FILL_25_DFFSR_49 ( );
FILL FILL_26_DFFSR_49 ( );
FILL FILL_27_DFFSR_49 ( );
FILL FILL_28_DFFSR_49 ( );
FILL FILL_29_DFFSR_49 ( );
FILL FILL_30_DFFSR_49 ( );
FILL FILL_31_DFFSR_49 ( );
FILL FILL_32_DFFSR_49 ( );
FILL FILL_33_DFFSR_49 ( );
FILL FILL_34_DFFSR_49 ( );
FILL FILL_35_DFFSR_49 ( );
FILL FILL_36_DFFSR_49 ( );
FILL FILL_37_DFFSR_49 ( );
FILL FILL_38_DFFSR_49 ( );
FILL FILL_39_DFFSR_49 ( );
FILL FILL_40_DFFSR_49 ( );
FILL FILL_41_DFFSR_49 ( );
FILL FILL_42_DFFSR_49 ( );
FILL FILL_43_DFFSR_49 ( );
FILL FILL_44_DFFSR_49 ( );
FILL FILL_45_DFFSR_49 ( );
FILL FILL_46_DFFSR_49 ( );
FILL FILL_47_DFFSR_49 ( );
FILL FILL_48_DFFSR_49 ( );
FILL FILL_49_DFFSR_49 ( );
FILL FILL_50_DFFSR_49 ( );
FILL FILL_0_CLKBUF1_40 ( );
FILL FILL_1_CLKBUF1_40 ( );
FILL FILL_2_CLKBUF1_40 ( );
FILL FILL_3_CLKBUF1_40 ( );
FILL FILL_4_CLKBUF1_40 ( );
FILL FILL_5_CLKBUF1_40 ( );
FILL FILL_6_CLKBUF1_40 ( );
FILL FILL_7_CLKBUF1_40 ( );
FILL FILL_8_CLKBUF1_40 ( );
FILL FILL_9_CLKBUF1_40 ( );
FILL FILL_10_CLKBUF1_40 ( );
FILL FILL_11_CLKBUF1_40 ( );
FILL FILL_12_CLKBUF1_40 ( );
FILL FILL_13_CLKBUF1_40 ( );
FILL FILL_14_CLKBUF1_40 ( );
FILL FILL_15_CLKBUF1_40 ( );
FILL FILL_16_CLKBUF1_40 ( );
FILL FILL_17_CLKBUF1_40 ( );
FILL FILL_18_CLKBUF1_40 ( );
FILL FILL_19_CLKBUF1_40 ( );
FILL FILL_20_CLKBUF1_40 ( );
FILL FILL_0_DFFSR_170 ( );
FILL FILL_1_DFFSR_170 ( );
FILL FILL_2_DFFSR_170 ( );
FILL FILL_3_DFFSR_170 ( );
FILL FILL_4_DFFSR_170 ( );
FILL FILL_5_DFFSR_170 ( );
FILL FILL_6_DFFSR_170 ( );
FILL FILL_7_DFFSR_170 ( );
FILL FILL_8_DFFSR_170 ( );
FILL FILL_9_DFFSR_170 ( );
FILL FILL_10_DFFSR_170 ( );
FILL FILL_11_DFFSR_170 ( );
FILL FILL_12_DFFSR_170 ( );
FILL FILL_13_DFFSR_170 ( );
FILL FILL_14_DFFSR_170 ( );
FILL FILL_15_DFFSR_170 ( );
FILL FILL_16_DFFSR_170 ( );
FILL FILL_17_DFFSR_170 ( );
FILL FILL_18_DFFSR_170 ( );
FILL FILL_19_DFFSR_170 ( );
FILL FILL_20_DFFSR_170 ( );
FILL FILL_21_DFFSR_170 ( );
FILL FILL_22_DFFSR_170 ( );
FILL FILL_23_DFFSR_170 ( );
FILL FILL_24_DFFSR_170 ( );
FILL FILL_25_DFFSR_170 ( );
FILL FILL_26_DFFSR_170 ( );
FILL FILL_27_DFFSR_170 ( );
FILL FILL_28_DFFSR_170 ( );
FILL FILL_29_DFFSR_170 ( );
FILL FILL_30_DFFSR_170 ( );
FILL FILL_31_DFFSR_170 ( );
FILL FILL_32_DFFSR_170 ( );
FILL FILL_33_DFFSR_170 ( );
FILL FILL_34_DFFSR_170 ( );
FILL FILL_35_DFFSR_170 ( );
FILL FILL_36_DFFSR_170 ( );
FILL FILL_37_DFFSR_170 ( );
FILL FILL_38_DFFSR_170 ( );
FILL FILL_39_DFFSR_170 ( );
FILL FILL_40_DFFSR_170 ( );
FILL FILL_41_DFFSR_170 ( );
FILL FILL_42_DFFSR_170 ( );
FILL FILL_43_DFFSR_170 ( );
FILL FILL_44_DFFSR_170 ( );
FILL FILL_45_DFFSR_170 ( );
FILL FILL_46_DFFSR_170 ( );
FILL FILL_47_DFFSR_170 ( );
FILL FILL_48_DFFSR_170 ( );
FILL FILL_49_DFFSR_170 ( );
FILL FILL_50_DFFSR_170 ( );
FILL FILL_51_DFFSR_170 ( );
FILL FILL_0_NOR2X1_39 ( );
FILL FILL_1_NOR2X1_39 ( );
FILL FILL_2_NOR2X1_39 ( );
FILL FILL_3_NOR2X1_39 ( );
FILL FILL_4_NOR2X1_39 ( );
FILL FILL_5_NOR2X1_39 ( );
FILL FILL_6_NOR2X1_39 ( );
FILL FILL_0_DFFSR_168 ( );
FILL FILL_1_DFFSR_168 ( );
FILL FILL_2_DFFSR_168 ( );
FILL FILL_3_DFFSR_168 ( );
FILL FILL_4_DFFSR_168 ( );
FILL FILL_5_DFFSR_168 ( );
FILL FILL_6_DFFSR_168 ( );
FILL FILL_7_DFFSR_168 ( );
FILL FILL_8_DFFSR_168 ( );
FILL FILL_9_DFFSR_168 ( );
FILL FILL_10_DFFSR_168 ( );
FILL FILL_11_DFFSR_168 ( );
FILL FILL_12_DFFSR_168 ( );
FILL FILL_13_DFFSR_168 ( );
FILL FILL_14_DFFSR_168 ( );
FILL FILL_15_DFFSR_168 ( );
FILL FILL_16_DFFSR_168 ( );
FILL FILL_17_DFFSR_168 ( );
FILL FILL_18_DFFSR_168 ( );
FILL FILL_19_DFFSR_168 ( );
FILL FILL_20_DFFSR_168 ( );
FILL FILL_21_DFFSR_168 ( );
FILL FILL_22_DFFSR_168 ( );
FILL FILL_23_DFFSR_168 ( );
FILL FILL_24_DFFSR_168 ( );
FILL FILL_25_DFFSR_168 ( );
FILL FILL_26_DFFSR_168 ( );
FILL FILL_27_DFFSR_168 ( );
FILL FILL_28_DFFSR_168 ( );
FILL FILL_29_DFFSR_168 ( );
FILL FILL_30_DFFSR_168 ( );
FILL FILL_31_DFFSR_168 ( );
FILL FILL_32_DFFSR_168 ( );
FILL FILL_33_DFFSR_168 ( );
FILL FILL_34_DFFSR_168 ( );
FILL FILL_35_DFFSR_168 ( );
FILL FILL_36_DFFSR_168 ( );
FILL FILL_37_DFFSR_168 ( );
FILL FILL_38_DFFSR_168 ( );
FILL FILL_39_DFFSR_168 ( );
FILL FILL_40_DFFSR_168 ( );
FILL FILL_41_DFFSR_168 ( );
FILL FILL_42_DFFSR_168 ( );
FILL FILL_43_DFFSR_168 ( );
FILL FILL_44_DFFSR_168 ( );
FILL FILL_45_DFFSR_168 ( );
FILL FILL_46_DFFSR_168 ( );
FILL FILL_47_DFFSR_168 ( );
FILL FILL_48_DFFSR_168 ( );
FILL FILL_49_DFFSR_168 ( );
FILL FILL_50_DFFSR_168 ( );
FILL FILL_0_INVX1_165 ( );
FILL FILL_1_INVX1_165 ( );
FILL FILL_2_INVX1_165 ( );
FILL FILL_3_INVX1_165 ( );
FILL FILL_4_INVX1_165 ( );
FILL FILL_0_DFFSR_275 ( );
FILL FILL_1_DFFSR_275 ( );
FILL FILL_2_DFFSR_275 ( );
FILL FILL_3_DFFSR_275 ( );
FILL FILL_4_DFFSR_275 ( );
FILL FILL_5_DFFSR_275 ( );
FILL FILL_6_DFFSR_275 ( );
FILL FILL_7_DFFSR_275 ( );
FILL FILL_8_DFFSR_275 ( );
FILL FILL_9_DFFSR_275 ( );
FILL FILL_10_DFFSR_275 ( );
FILL FILL_11_DFFSR_275 ( );
FILL FILL_12_DFFSR_275 ( );
FILL FILL_13_DFFSR_275 ( );
FILL FILL_14_DFFSR_275 ( );
FILL FILL_15_DFFSR_275 ( );
FILL FILL_16_DFFSR_275 ( );
FILL FILL_17_DFFSR_275 ( );
FILL FILL_18_DFFSR_275 ( );
FILL FILL_19_DFFSR_275 ( );
FILL FILL_20_DFFSR_275 ( );
FILL FILL_21_DFFSR_275 ( );
FILL FILL_22_DFFSR_275 ( );
FILL FILL_23_DFFSR_275 ( );
FILL FILL_24_DFFSR_275 ( );
FILL FILL_25_DFFSR_275 ( );
FILL FILL_26_DFFSR_275 ( );
FILL FILL_27_DFFSR_275 ( );
FILL FILL_28_DFFSR_275 ( );
FILL FILL_29_DFFSR_275 ( );
FILL FILL_30_DFFSR_275 ( );
FILL FILL_31_DFFSR_275 ( );
FILL FILL_32_DFFSR_275 ( );
FILL FILL_33_DFFSR_275 ( );
FILL FILL_34_DFFSR_275 ( );
FILL FILL_35_DFFSR_275 ( );
FILL FILL_36_DFFSR_275 ( );
FILL FILL_37_DFFSR_275 ( );
FILL FILL_38_DFFSR_275 ( );
FILL FILL_39_DFFSR_275 ( );
FILL FILL_40_DFFSR_275 ( );
FILL FILL_41_DFFSR_275 ( );
FILL FILL_42_DFFSR_275 ( );
FILL FILL_43_DFFSR_275 ( );
FILL FILL_44_DFFSR_275 ( );
FILL FILL_45_DFFSR_275 ( );
FILL FILL_46_DFFSR_275 ( );
FILL FILL_47_DFFSR_275 ( );
FILL FILL_48_DFFSR_275 ( );
FILL FILL_49_DFFSR_275 ( );
FILL FILL_50_DFFSR_275 ( );
FILL FILL_51_DFFSR_275 ( );
FILL FILL_0_DFFPOSX1_49 ( );
FILL FILL_1_DFFPOSX1_49 ( );
FILL FILL_2_DFFPOSX1_49 ( );
FILL FILL_3_DFFPOSX1_49 ( );
FILL FILL_4_DFFPOSX1_49 ( );
FILL FILL_5_DFFPOSX1_49 ( );
FILL FILL_6_DFFPOSX1_49 ( );
FILL FILL_7_DFFPOSX1_49 ( );
FILL FILL_8_DFFPOSX1_49 ( );
FILL FILL_9_DFFPOSX1_49 ( );
FILL FILL_10_DFFPOSX1_49 ( );
FILL FILL_11_DFFPOSX1_49 ( );
FILL FILL_12_DFFPOSX1_49 ( );
FILL FILL_13_DFFPOSX1_49 ( );
FILL FILL_14_DFFPOSX1_49 ( );
FILL FILL_15_DFFPOSX1_49 ( );
FILL FILL_16_DFFPOSX1_49 ( );
FILL FILL_17_DFFPOSX1_49 ( );
FILL FILL_18_DFFPOSX1_49 ( );
FILL FILL_19_DFFPOSX1_49 ( );
FILL FILL_20_DFFPOSX1_49 ( );
FILL FILL_21_DFFPOSX1_49 ( );
FILL FILL_22_DFFPOSX1_49 ( );
FILL FILL_23_DFFPOSX1_49 ( );
FILL FILL_24_DFFPOSX1_49 ( );
FILL FILL_25_DFFPOSX1_49 ( );
FILL FILL_26_DFFPOSX1_49 ( );
FILL FILL_27_DFFPOSX1_49 ( );
FILL FILL_0_INVX1_205 ( );
FILL FILL_1_INVX1_205 ( );
FILL FILL_2_INVX1_205 ( );
FILL FILL_3_INVX1_205 ( );
FILL FILL_4_INVX1_205 ( );
FILL FILL_0_DFFSR_92 ( );
FILL FILL_1_DFFSR_92 ( );
FILL FILL_2_DFFSR_92 ( );
FILL FILL_3_DFFSR_92 ( );
FILL FILL_4_DFFSR_92 ( );
FILL FILL_5_DFFSR_92 ( );
FILL FILL_6_DFFSR_92 ( );
FILL FILL_7_DFFSR_92 ( );
FILL FILL_8_DFFSR_92 ( );
FILL FILL_9_DFFSR_92 ( );
FILL FILL_10_DFFSR_92 ( );
FILL FILL_11_DFFSR_92 ( );
FILL FILL_12_DFFSR_92 ( );
FILL FILL_13_DFFSR_92 ( );
FILL FILL_14_DFFSR_92 ( );
FILL FILL_15_DFFSR_92 ( );
FILL FILL_16_DFFSR_92 ( );
FILL FILL_17_DFFSR_92 ( );
FILL FILL_18_DFFSR_92 ( );
FILL FILL_19_DFFSR_92 ( );
FILL FILL_20_DFFSR_92 ( );
FILL FILL_21_DFFSR_92 ( );
FILL FILL_22_DFFSR_92 ( );
FILL FILL_23_DFFSR_92 ( );
FILL FILL_24_DFFSR_92 ( );
FILL FILL_25_DFFSR_92 ( );
FILL FILL_26_DFFSR_92 ( );
FILL FILL_27_DFFSR_92 ( );
FILL FILL_28_DFFSR_92 ( );
FILL FILL_29_DFFSR_92 ( );
FILL FILL_30_DFFSR_92 ( );
FILL FILL_31_DFFSR_92 ( );
FILL FILL_32_DFFSR_92 ( );
FILL FILL_33_DFFSR_92 ( );
FILL FILL_34_DFFSR_92 ( );
FILL FILL_35_DFFSR_92 ( );
FILL FILL_36_DFFSR_92 ( );
FILL FILL_37_DFFSR_92 ( );
FILL FILL_38_DFFSR_92 ( );
FILL FILL_39_DFFSR_92 ( );
FILL FILL_40_DFFSR_92 ( );
FILL FILL_41_DFFSR_92 ( );
FILL FILL_42_DFFSR_92 ( );
FILL FILL_43_DFFSR_92 ( );
FILL FILL_44_DFFSR_92 ( );
FILL FILL_45_DFFSR_92 ( );
FILL FILL_46_DFFSR_92 ( );
FILL FILL_47_DFFSR_92 ( );
FILL FILL_48_DFFSR_92 ( );
FILL FILL_49_DFFSR_92 ( );
FILL FILL_50_DFFSR_92 ( );
FILL FILL_51_DFFSR_92 ( );
FILL FILL_0_AOI22X1_4 ( );
FILL FILL_1_AOI22X1_4 ( );
FILL FILL_2_AOI22X1_4 ( );
FILL FILL_3_AOI22X1_4 ( );
FILL FILL_4_AOI22X1_4 ( );
FILL FILL_5_AOI22X1_4 ( );
FILL FILL_6_AOI22X1_4 ( );
FILL FILL_7_AOI22X1_4 ( );
FILL FILL_8_AOI22X1_4 ( );
FILL FILL_9_AOI22X1_4 ( );
FILL FILL_10_AOI22X1_4 ( );
FILL FILL_11_AOI22X1_4 ( );
FILL FILL_0_OAI22X1_11 ( );
FILL FILL_1_OAI22X1_11 ( );
FILL FILL_2_OAI22X1_11 ( );
FILL FILL_3_OAI22X1_11 ( );
FILL FILL_4_OAI22X1_11 ( );
FILL FILL_5_OAI22X1_11 ( );
FILL FILL_6_OAI22X1_11 ( );
FILL FILL_7_OAI22X1_11 ( );
FILL FILL_8_OAI22X1_11 ( );
FILL FILL_9_OAI22X1_11 ( );
FILL FILL_10_OAI22X1_11 ( );
FILL FILL_11_OAI22X1_11 ( );
FILL FILL_0_NOR2X1_1 ( );
FILL FILL_1_NOR2X1_1 ( );
FILL FILL_2_NOR2X1_1 ( );
FILL FILL_3_NOR2X1_1 ( );
FILL FILL_4_NOR2X1_1 ( );
FILL FILL_5_NOR2X1_1 ( );
FILL FILL_6_NOR2X1_1 ( );
FILL FILL_0_AOI21X1_71 ( );
FILL FILL_1_AOI21X1_71 ( );
FILL FILL_2_AOI21X1_71 ( );
FILL FILL_3_AOI21X1_71 ( );
FILL FILL_4_AOI21X1_71 ( );
FILL FILL_5_AOI21X1_71 ( );
FILL FILL_6_AOI21X1_71 ( );
FILL FILL_7_AOI21X1_71 ( );
FILL FILL_8_AOI21X1_71 ( );
FILL FILL_9_AOI21X1_71 ( );
FILL FILL_0_NAND2X1_181 ( );
FILL FILL_1_NAND2X1_181 ( );
FILL FILL_2_NAND2X1_181 ( );
FILL FILL_3_NAND2X1_181 ( );
FILL FILL_4_NAND2X1_181 ( );
FILL FILL_5_NAND2X1_181 ( );
FILL FILL_6_NAND2X1_181 ( );
FILL FILL_0_DFFSR_127 ( );
FILL FILL_1_DFFSR_127 ( );
FILL FILL_2_DFFSR_127 ( );
FILL FILL_3_DFFSR_127 ( );
FILL FILL_4_DFFSR_127 ( );
FILL FILL_5_DFFSR_127 ( );
FILL FILL_6_DFFSR_127 ( );
FILL FILL_7_DFFSR_127 ( );
FILL FILL_8_DFFSR_127 ( );
FILL FILL_9_DFFSR_127 ( );
FILL FILL_10_DFFSR_127 ( );
FILL FILL_11_DFFSR_127 ( );
FILL FILL_12_DFFSR_127 ( );
FILL FILL_13_DFFSR_127 ( );
FILL FILL_14_DFFSR_127 ( );
FILL FILL_15_DFFSR_127 ( );
FILL FILL_16_DFFSR_127 ( );
FILL FILL_17_DFFSR_127 ( );
FILL FILL_18_DFFSR_127 ( );
FILL FILL_19_DFFSR_127 ( );
FILL FILL_20_DFFSR_127 ( );
FILL FILL_21_DFFSR_127 ( );
FILL FILL_22_DFFSR_127 ( );
FILL FILL_23_DFFSR_127 ( );
FILL FILL_24_DFFSR_127 ( );
FILL FILL_25_DFFSR_127 ( );
FILL FILL_26_DFFSR_127 ( );
FILL FILL_27_DFFSR_127 ( );
FILL FILL_28_DFFSR_127 ( );
FILL FILL_29_DFFSR_127 ( );
FILL FILL_30_DFFSR_127 ( );
FILL FILL_31_DFFSR_127 ( );
FILL FILL_32_DFFSR_127 ( );
FILL FILL_33_DFFSR_127 ( );
FILL FILL_34_DFFSR_127 ( );
FILL FILL_35_DFFSR_127 ( );
FILL FILL_36_DFFSR_127 ( );
FILL FILL_37_DFFSR_127 ( );
FILL FILL_38_DFFSR_127 ( );
FILL FILL_39_DFFSR_127 ( );
FILL FILL_40_DFFSR_127 ( );
FILL FILL_41_DFFSR_127 ( );
FILL FILL_42_DFFSR_127 ( );
FILL FILL_43_DFFSR_127 ( );
FILL FILL_44_DFFSR_127 ( );
FILL FILL_45_DFFSR_127 ( );
FILL FILL_46_DFFSR_127 ( );
FILL FILL_47_DFFSR_127 ( );
FILL FILL_48_DFFSR_127 ( );
FILL FILL_49_DFFSR_127 ( );
FILL FILL_50_DFFSR_127 ( );
FILL FILL_0_CLKBUF1_5 ( );
FILL FILL_1_CLKBUF1_5 ( );
FILL FILL_2_CLKBUF1_5 ( );
FILL FILL_3_CLKBUF1_5 ( );
FILL FILL_4_CLKBUF1_5 ( );
FILL FILL_5_CLKBUF1_5 ( );
FILL FILL_6_CLKBUF1_5 ( );
FILL FILL_7_CLKBUF1_5 ( );
FILL FILL_8_CLKBUF1_5 ( );
FILL FILL_9_CLKBUF1_5 ( );
FILL FILL_10_CLKBUF1_5 ( );
FILL FILL_11_CLKBUF1_5 ( );
FILL FILL_12_CLKBUF1_5 ( );
FILL FILL_13_CLKBUF1_5 ( );
FILL FILL_14_CLKBUF1_5 ( );
FILL FILL_15_CLKBUF1_5 ( );
FILL FILL_16_CLKBUF1_5 ( );
FILL FILL_17_CLKBUF1_5 ( );
FILL FILL_18_CLKBUF1_5 ( );
FILL FILL_19_CLKBUF1_5 ( );
FILL FILL_20_CLKBUF1_5 ( );
FILL FILL_0_NAND3X1_6 ( );
FILL FILL_1_NAND3X1_6 ( );
FILL FILL_2_NAND3X1_6 ( );
FILL FILL_3_NAND3X1_6 ( );
FILL FILL_4_NAND3X1_6 ( );
FILL FILL_5_NAND3X1_6 ( );
FILL FILL_6_NAND3X1_6 ( );
FILL FILL_7_NAND3X1_6 ( );
FILL FILL_8_NAND3X1_6 ( );
FILL FILL_9_NAND3X1_6 ( );
FILL FILL_0_NOR2X1_13 ( );
FILL FILL_1_NOR2X1_13 ( );
FILL FILL_2_NOR2X1_13 ( );
FILL FILL_3_NOR2X1_13 ( );
FILL FILL_4_NOR2X1_13 ( );
FILL FILL_5_NOR2X1_13 ( );
FILL FILL_6_NOR2X1_13 ( );
FILL FILL_0_NAND2X1_15 ( );
FILL FILL_1_NAND2X1_15 ( );
FILL FILL_2_NAND2X1_15 ( );
FILL FILL_3_NAND2X1_15 ( );
FILL FILL_4_NAND2X1_15 ( );
FILL FILL_5_NAND2X1_15 ( );
FILL FILL_6_NAND2X1_15 ( );
FILL FILL_0_OAI21X1_3 ( );
FILL FILL_1_OAI21X1_3 ( );
FILL FILL_2_OAI21X1_3 ( );
FILL FILL_3_OAI21X1_3 ( );
FILL FILL_4_OAI21X1_3 ( );
FILL FILL_5_OAI21X1_3 ( );
FILL FILL_6_OAI21X1_3 ( );
FILL FILL_7_OAI21X1_3 ( );
FILL FILL_8_OAI21X1_3 ( );
FILL FILL_0_NAND3X1_19 ( );
FILL FILL_1_NAND3X1_19 ( );
FILL FILL_2_NAND3X1_19 ( );
FILL FILL_3_NAND3X1_19 ( );
FILL FILL_4_NAND3X1_19 ( );
FILL FILL_5_NAND3X1_19 ( );
FILL FILL_6_NAND3X1_19 ( );
FILL FILL_7_NAND3X1_19 ( );
FILL FILL_8_NAND3X1_19 ( );
FILL FILL_0_NAND3X1_3 ( );
FILL FILL_1_NAND3X1_3 ( );
FILL FILL_2_NAND3X1_3 ( );
FILL FILL_3_NAND3X1_3 ( );
FILL FILL_4_NAND3X1_3 ( );
FILL FILL_5_NAND3X1_3 ( );
FILL FILL_6_NAND3X1_3 ( );
FILL FILL_7_NAND3X1_3 ( );
FILL FILL_8_NAND3X1_3 ( );
FILL FILL_0_NAND2X1_13 ( );
FILL FILL_1_NAND2X1_13 ( );
FILL FILL_2_NAND2X1_13 ( );
FILL FILL_3_NAND2X1_13 ( );
FILL FILL_4_NAND2X1_13 ( );
FILL FILL_5_NAND2X1_13 ( );
FILL FILL_6_NAND2X1_13 ( );
FILL FILL_0_DFFSR_113 ( );
FILL FILL_1_DFFSR_113 ( );
FILL FILL_2_DFFSR_113 ( );
FILL FILL_3_DFFSR_113 ( );
FILL FILL_4_DFFSR_113 ( );
FILL FILL_5_DFFSR_113 ( );
FILL FILL_6_DFFSR_113 ( );
FILL FILL_7_DFFSR_113 ( );
FILL FILL_8_DFFSR_113 ( );
FILL FILL_9_DFFSR_113 ( );
FILL FILL_10_DFFSR_113 ( );
FILL FILL_11_DFFSR_113 ( );
FILL FILL_12_DFFSR_113 ( );
FILL FILL_13_DFFSR_113 ( );
FILL FILL_14_DFFSR_113 ( );
FILL FILL_15_DFFSR_113 ( );
FILL FILL_16_DFFSR_113 ( );
FILL FILL_17_DFFSR_113 ( );
FILL FILL_18_DFFSR_113 ( );
FILL FILL_19_DFFSR_113 ( );
FILL FILL_20_DFFSR_113 ( );
FILL FILL_21_DFFSR_113 ( );
FILL FILL_22_DFFSR_113 ( );
FILL FILL_23_DFFSR_113 ( );
FILL FILL_24_DFFSR_113 ( );
FILL FILL_25_DFFSR_113 ( );
FILL FILL_26_DFFSR_113 ( );
FILL FILL_27_DFFSR_113 ( );
FILL FILL_28_DFFSR_113 ( );
FILL FILL_29_DFFSR_113 ( );
FILL FILL_30_DFFSR_113 ( );
FILL FILL_31_DFFSR_113 ( );
FILL FILL_32_DFFSR_113 ( );
FILL FILL_33_DFFSR_113 ( );
FILL FILL_34_DFFSR_113 ( );
FILL FILL_35_DFFSR_113 ( );
FILL FILL_36_DFFSR_113 ( );
FILL FILL_37_DFFSR_113 ( );
FILL FILL_38_DFFSR_113 ( );
FILL FILL_39_DFFSR_113 ( );
FILL FILL_40_DFFSR_113 ( );
FILL FILL_41_DFFSR_113 ( );
FILL FILL_42_DFFSR_113 ( );
FILL FILL_43_DFFSR_113 ( );
FILL FILL_44_DFFSR_113 ( );
FILL FILL_45_DFFSR_113 ( );
FILL FILL_46_DFFSR_113 ( );
FILL FILL_47_DFFSR_113 ( );
FILL FILL_48_DFFSR_113 ( );
FILL FILL_49_DFFSR_113 ( );
FILL FILL_50_DFFSR_113 ( );
FILL FILL_0_DFFSR_162 ( );
FILL FILL_1_DFFSR_162 ( );
FILL FILL_2_DFFSR_162 ( );
FILL FILL_3_DFFSR_162 ( );
FILL FILL_4_DFFSR_162 ( );
FILL FILL_5_DFFSR_162 ( );
FILL FILL_6_DFFSR_162 ( );
FILL FILL_7_DFFSR_162 ( );
FILL FILL_8_DFFSR_162 ( );
FILL FILL_9_DFFSR_162 ( );
FILL FILL_10_DFFSR_162 ( );
FILL FILL_11_DFFSR_162 ( );
FILL FILL_12_DFFSR_162 ( );
FILL FILL_13_DFFSR_162 ( );
FILL FILL_14_DFFSR_162 ( );
FILL FILL_15_DFFSR_162 ( );
FILL FILL_16_DFFSR_162 ( );
FILL FILL_17_DFFSR_162 ( );
FILL FILL_18_DFFSR_162 ( );
FILL FILL_19_DFFSR_162 ( );
FILL FILL_20_DFFSR_162 ( );
FILL FILL_21_DFFSR_162 ( );
FILL FILL_22_DFFSR_162 ( );
FILL FILL_23_DFFSR_162 ( );
FILL FILL_24_DFFSR_162 ( );
FILL FILL_25_DFFSR_162 ( );
FILL FILL_26_DFFSR_162 ( );
FILL FILL_27_DFFSR_162 ( );
FILL FILL_28_DFFSR_162 ( );
FILL FILL_29_DFFSR_162 ( );
FILL FILL_30_DFFSR_162 ( );
FILL FILL_31_DFFSR_162 ( );
FILL FILL_32_DFFSR_162 ( );
FILL FILL_33_DFFSR_162 ( );
FILL FILL_34_DFFSR_162 ( );
FILL FILL_35_DFFSR_162 ( );
FILL FILL_36_DFFSR_162 ( );
FILL FILL_37_DFFSR_162 ( );
FILL FILL_38_DFFSR_162 ( );
FILL FILL_39_DFFSR_162 ( );
FILL FILL_40_DFFSR_162 ( );
FILL FILL_41_DFFSR_162 ( );
FILL FILL_42_DFFSR_162 ( );
FILL FILL_43_DFFSR_162 ( );
FILL FILL_44_DFFSR_162 ( );
FILL FILL_45_DFFSR_162 ( );
FILL FILL_46_DFFSR_162 ( );
FILL FILL_47_DFFSR_162 ( );
FILL FILL_48_DFFSR_162 ( );
FILL FILL_49_DFFSR_162 ( );
FILL FILL_50_DFFSR_162 ( );
FILL FILL_0_INVX1_74 ( );
FILL FILL_1_INVX1_74 ( );
FILL FILL_2_INVX1_74 ( );
FILL FILL_3_INVX1_74 ( );
FILL FILL_4_INVX1_74 ( );
FILL FILL_0_DFFSR_186 ( );
FILL FILL_1_DFFSR_186 ( );
FILL FILL_2_DFFSR_186 ( );
FILL FILL_3_DFFSR_186 ( );
FILL FILL_4_DFFSR_186 ( );
FILL FILL_5_DFFSR_186 ( );
FILL FILL_6_DFFSR_186 ( );
FILL FILL_7_DFFSR_186 ( );
FILL FILL_8_DFFSR_186 ( );
FILL FILL_9_DFFSR_186 ( );
FILL FILL_10_DFFSR_186 ( );
FILL FILL_11_DFFSR_186 ( );
FILL FILL_12_DFFSR_186 ( );
FILL FILL_13_DFFSR_186 ( );
FILL FILL_14_DFFSR_186 ( );
FILL FILL_15_DFFSR_186 ( );
FILL FILL_16_DFFSR_186 ( );
FILL FILL_17_DFFSR_186 ( );
FILL FILL_18_DFFSR_186 ( );
FILL FILL_19_DFFSR_186 ( );
FILL FILL_20_DFFSR_186 ( );
FILL FILL_21_DFFSR_186 ( );
FILL FILL_22_DFFSR_186 ( );
FILL FILL_23_DFFSR_186 ( );
FILL FILL_24_DFFSR_186 ( );
FILL FILL_25_DFFSR_186 ( );
FILL FILL_26_DFFSR_186 ( );
FILL FILL_27_DFFSR_186 ( );
FILL FILL_28_DFFSR_186 ( );
FILL FILL_29_DFFSR_186 ( );
FILL FILL_30_DFFSR_186 ( );
FILL FILL_31_DFFSR_186 ( );
FILL FILL_32_DFFSR_186 ( );
FILL FILL_33_DFFSR_186 ( );
FILL FILL_34_DFFSR_186 ( );
FILL FILL_35_DFFSR_186 ( );
FILL FILL_36_DFFSR_186 ( );
FILL FILL_37_DFFSR_186 ( );
FILL FILL_38_DFFSR_186 ( );
FILL FILL_39_DFFSR_186 ( );
FILL FILL_40_DFFSR_186 ( );
FILL FILL_41_DFFSR_186 ( );
FILL FILL_42_DFFSR_186 ( );
FILL FILL_43_DFFSR_186 ( );
FILL FILL_44_DFFSR_186 ( );
FILL FILL_45_DFFSR_186 ( );
FILL FILL_46_DFFSR_186 ( );
FILL FILL_47_DFFSR_186 ( );
FILL FILL_48_DFFSR_186 ( );
FILL FILL_49_DFFSR_186 ( );
FILL FILL_50_DFFSR_186 ( );
FILL FILL_0_XOR2X1_6 ( );
FILL FILL_1_XOR2X1_6 ( );
FILL FILL_2_XOR2X1_6 ( );
FILL FILL_3_XOR2X1_6 ( );
FILL FILL_4_XOR2X1_6 ( );
FILL FILL_5_XOR2X1_6 ( );
FILL FILL_6_XOR2X1_6 ( );
FILL FILL_7_XOR2X1_6 ( );
FILL FILL_8_XOR2X1_6 ( );
FILL FILL_9_XOR2X1_6 ( );
FILL FILL_10_XOR2X1_6 ( );
FILL FILL_11_XOR2X1_6 ( );
FILL FILL_12_XOR2X1_6 ( );
FILL FILL_13_XOR2X1_6 ( );
FILL FILL_14_XOR2X1_6 ( );
FILL FILL_15_XOR2X1_6 ( );
FILL FILL_16_XOR2X1_6 ( );
FILL FILL_0_BUFX2_99 ( );
FILL FILL_1_BUFX2_99 ( );
FILL FILL_2_BUFX2_99 ( );
FILL FILL_3_BUFX2_99 ( );
FILL FILL_4_BUFX2_99 ( );
FILL FILL_5_BUFX2_99 ( );
FILL FILL_6_BUFX2_99 ( );
FILL FILL_0_INVX1_175 ( );
FILL FILL_1_INVX1_175 ( );
FILL FILL_2_INVX1_175 ( );
FILL FILL_3_INVX1_175 ( );
FILL FILL_4_INVX1_175 ( );
FILL FILL_0_DFFSR_279 ( );
FILL FILL_1_DFFSR_279 ( );
FILL FILL_2_DFFSR_279 ( );
FILL FILL_3_DFFSR_279 ( );
FILL FILL_4_DFFSR_279 ( );
FILL FILL_5_DFFSR_279 ( );
FILL FILL_6_DFFSR_279 ( );
FILL FILL_7_DFFSR_279 ( );
FILL FILL_8_DFFSR_279 ( );
FILL FILL_9_DFFSR_279 ( );
FILL FILL_10_DFFSR_279 ( );
FILL FILL_11_DFFSR_279 ( );
FILL FILL_12_DFFSR_279 ( );
FILL FILL_13_DFFSR_279 ( );
FILL FILL_14_DFFSR_279 ( );
FILL FILL_15_DFFSR_279 ( );
FILL FILL_16_DFFSR_279 ( );
FILL FILL_17_DFFSR_279 ( );
FILL FILL_18_DFFSR_279 ( );
FILL FILL_19_DFFSR_279 ( );
FILL FILL_20_DFFSR_279 ( );
FILL FILL_21_DFFSR_279 ( );
FILL FILL_22_DFFSR_279 ( );
FILL FILL_23_DFFSR_279 ( );
FILL FILL_24_DFFSR_279 ( );
FILL FILL_25_DFFSR_279 ( );
FILL FILL_26_DFFSR_279 ( );
FILL FILL_27_DFFSR_279 ( );
FILL FILL_28_DFFSR_279 ( );
FILL FILL_29_DFFSR_279 ( );
FILL FILL_30_DFFSR_279 ( );
FILL FILL_31_DFFSR_279 ( );
FILL FILL_32_DFFSR_279 ( );
FILL FILL_33_DFFSR_279 ( );
FILL FILL_34_DFFSR_279 ( );
FILL FILL_35_DFFSR_279 ( );
FILL FILL_36_DFFSR_279 ( );
FILL FILL_37_DFFSR_279 ( );
FILL FILL_38_DFFSR_279 ( );
FILL FILL_39_DFFSR_279 ( );
FILL FILL_40_DFFSR_279 ( );
FILL FILL_41_DFFSR_279 ( );
FILL FILL_42_DFFSR_279 ( );
FILL FILL_43_DFFSR_279 ( );
FILL FILL_44_DFFSR_279 ( );
FILL FILL_45_DFFSR_279 ( );
FILL FILL_46_DFFSR_279 ( );
FILL FILL_47_DFFSR_279 ( );
FILL FILL_48_DFFSR_279 ( );
FILL FILL_49_DFFSR_279 ( );
FILL FILL_50_DFFSR_279 ( );
FILL FILL_0_DFFSR_84 ( );
FILL FILL_1_DFFSR_84 ( );
FILL FILL_2_DFFSR_84 ( );
FILL FILL_3_DFFSR_84 ( );
FILL FILL_4_DFFSR_84 ( );
FILL FILL_5_DFFSR_84 ( );
FILL FILL_6_DFFSR_84 ( );
FILL FILL_7_DFFSR_84 ( );
FILL FILL_8_DFFSR_84 ( );
FILL FILL_9_DFFSR_84 ( );
FILL FILL_10_DFFSR_84 ( );
FILL FILL_11_DFFSR_84 ( );
FILL FILL_12_DFFSR_84 ( );
FILL FILL_13_DFFSR_84 ( );
FILL FILL_14_DFFSR_84 ( );
FILL FILL_15_DFFSR_84 ( );
FILL FILL_16_DFFSR_84 ( );
FILL FILL_17_DFFSR_84 ( );
FILL FILL_18_DFFSR_84 ( );
FILL FILL_19_DFFSR_84 ( );
FILL FILL_20_DFFSR_84 ( );
FILL FILL_21_DFFSR_84 ( );
FILL FILL_22_DFFSR_84 ( );
FILL FILL_23_DFFSR_84 ( );
FILL FILL_24_DFFSR_84 ( );
FILL FILL_25_DFFSR_84 ( );
FILL FILL_26_DFFSR_84 ( );
FILL FILL_27_DFFSR_84 ( );
FILL FILL_28_DFFSR_84 ( );
FILL FILL_29_DFFSR_84 ( );
FILL FILL_30_DFFSR_84 ( );
FILL FILL_31_DFFSR_84 ( );
FILL FILL_32_DFFSR_84 ( );
FILL FILL_33_DFFSR_84 ( );
FILL FILL_34_DFFSR_84 ( );
FILL FILL_35_DFFSR_84 ( );
FILL FILL_36_DFFSR_84 ( );
FILL FILL_37_DFFSR_84 ( );
FILL FILL_38_DFFSR_84 ( );
FILL FILL_39_DFFSR_84 ( );
FILL FILL_40_DFFSR_84 ( );
FILL FILL_41_DFFSR_84 ( );
FILL FILL_42_DFFSR_84 ( );
FILL FILL_43_DFFSR_84 ( );
FILL FILL_44_DFFSR_84 ( );
FILL FILL_45_DFFSR_84 ( );
FILL FILL_46_DFFSR_84 ( );
FILL FILL_47_DFFSR_84 ( );
FILL FILL_48_DFFSR_84 ( );
FILL FILL_49_DFFSR_84 ( );
FILL FILL_50_DFFSR_84 ( );
FILL FILL_0_INVX1_27 ( );
FILL FILL_1_INVX1_27 ( );
FILL FILL_2_INVX1_27 ( );
FILL FILL_3_INVX1_27 ( );
FILL FILL_4_INVX1_27 ( );
FILL FILL_0_INVX1_4 ( );
FILL FILL_1_INVX1_4 ( );
FILL FILL_2_INVX1_4 ( );
FILL FILL_3_INVX1_4 ( );
FILL FILL_0_AND2X2_2 ( );
FILL FILL_1_AND2X2_2 ( );
FILL FILL_2_AND2X2_2 ( );
FILL FILL_3_AND2X2_2 ( );
FILL FILL_4_AND2X2_2 ( );
FILL FILL_5_AND2X2_2 ( );
FILL FILL_6_AND2X2_2 ( );
FILL FILL_7_AND2X2_2 ( );
FILL FILL_8_AND2X2_2 ( );
FILL FILL_9_AND2X2_2 ( );
FILL FILL_0_NAND2X1_3 ( );
FILL FILL_1_NAND2X1_3 ( );
FILL FILL_2_NAND2X1_3 ( );
FILL FILL_3_NAND2X1_3 ( );
FILL FILL_4_NAND2X1_3 ( );
FILL FILL_5_NAND2X1_3 ( );
FILL FILL_6_NAND2X1_3 ( );
FILL FILL_0_NOR2X1_15 ( );
FILL FILL_1_NOR2X1_15 ( );
FILL FILL_2_NOR2X1_15 ( );
FILL FILL_3_NOR2X1_15 ( );
FILL FILL_4_NOR2X1_15 ( );
FILL FILL_5_NOR2X1_15 ( );
FILL FILL_6_NOR2X1_15 ( );
FILL FILL_0_NAND2X1_22 ( );
FILL FILL_1_NAND2X1_22 ( );
FILL FILL_2_NAND2X1_22 ( );
FILL FILL_3_NAND2X1_22 ( );
FILL FILL_4_NAND2X1_22 ( );
FILL FILL_5_NAND2X1_22 ( );
FILL FILL_6_NAND2X1_22 ( );
FILL FILL_0_XOR2X1_15 ( );
FILL FILL_1_XOR2X1_15 ( );
FILL FILL_2_XOR2X1_15 ( );
FILL FILL_3_XOR2X1_15 ( );
FILL FILL_4_XOR2X1_15 ( );
FILL FILL_5_XOR2X1_15 ( );
FILL FILL_6_XOR2X1_15 ( );
FILL FILL_7_XOR2X1_15 ( );
FILL FILL_8_XOR2X1_15 ( );
FILL FILL_9_XOR2X1_15 ( );
FILL FILL_10_XOR2X1_15 ( );
FILL FILL_11_XOR2X1_15 ( );
FILL FILL_12_XOR2X1_15 ( );
FILL FILL_13_XOR2X1_15 ( );
FILL FILL_14_XOR2X1_15 ( );
FILL FILL_15_XOR2X1_15 ( );
FILL FILL_0_NAND3X1_44 ( );
FILL FILL_1_NAND3X1_44 ( );
FILL FILL_2_NAND3X1_44 ( );
FILL FILL_3_NAND3X1_44 ( );
FILL FILL_4_NAND3X1_44 ( );
FILL FILL_5_NAND3X1_44 ( );
FILL FILL_6_NAND3X1_44 ( );
FILL FILL_7_NAND3X1_44 ( );
FILL FILL_8_NAND3X1_44 ( );
FILL FILL_9_NAND3X1_44 ( );
FILL FILL_0_AND2X2_11 ( );
FILL FILL_1_AND2X2_11 ( );
FILL FILL_2_AND2X2_11 ( );
FILL FILL_3_AND2X2_11 ( );
FILL FILL_4_AND2X2_11 ( );
FILL FILL_5_AND2X2_11 ( );
FILL FILL_6_AND2X2_11 ( );
FILL FILL_7_AND2X2_11 ( );
FILL FILL_8_AND2X2_11 ( );
FILL FILL_0_NAND2X1_2 ( );
FILL FILL_1_NAND2X1_2 ( );
FILL FILL_2_NAND2X1_2 ( );
FILL FILL_3_NAND2X1_2 ( );
FILL FILL_4_NAND2X1_2 ( );
FILL FILL_5_NAND2X1_2 ( );
FILL FILL_6_NAND2X1_2 ( );
FILL FILL_0_NAND3X1_51 ( );
FILL FILL_1_NAND3X1_51 ( );
FILL FILL_2_NAND3X1_51 ( );
FILL FILL_3_NAND3X1_51 ( );
FILL FILL_4_NAND3X1_51 ( );
FILL FILL_5_NAND3X1_51 ( );
FILL FILL_6_NAND3X1_51 ( );
FILL FILL_7_NAND3X1_51 ( );
FILL FILL_8_NAND3X1_51 ( );
FILL FILL_9_NAND3X1_51 ( );
FILL FILL_0_NAND3X1_43 ( );
FILL FILL_1_NAND3X1_43 ( );
FILL FILL_2_NAND3X1_43 ( );
FILL FILL_3_NAND3X1_43 ( );
FILL FILL_4_NAND3X1_43 ( );
FILL FILL_5_NAND3X1_43 ( );
FILL FILL_6_NAND3X1_43 ( );
FILL FILL_7_NAND3X1_43 ( );
FILL FILL_8_NAND3X1_43 ( );
FILL FILL_0_OAI21X1_8 ( );
FILL FILL_1_OAI21X1_8 ( );
FILL FILL_2_OAI21X1_8 ( );
FILL FILL_3_OAI21X1_8 ( );
FILL FILL_4_OAI21X1_8 ( );
FILL FILL_5_OAI21X1_8 ( );
FILL FILL_6_OAI21X1_8 ( );
FILL FILL_7_OAI21X1_8 ( );
FILL FILL_8_OAI21X1_8 ( );
FILL FILL_0_NAND2X1_25 ( );
FILL FILL_1_NAND2X1_25 ( );
FILL FILL_2_NAND2X1_25 ( );
FILL FILL_3_NAND2X1_25 ( );
FILL FILL_4_NAND2X1_25 ( );
FILL FILL_5_NAND2X1_25 ( );
FILL FILL_6_NAND2X1_25 ( );
FILL FILL_0_NAND3X1_5 ( );
FILL FILL_1_NAND3X1_5 ( );
FILL FILL_2_NAND3X1_5 ( );
FILL FILL_3_NAND3X1_5 ( );
FILL FILL_4_NAND3X1_5 ( );
FILL FILL_5_NAND3X1_5 ( );
FILL FILL_6_NAND3X1_5 ( );
FILL FILL_7_NAND3X1_5 ( );
FILL FILL_8_NAND3X1_5 ( );
FILL FILL_0_NAND3X1_17 ( );
FILL FILL_1_NAND3X1_17 ( );
FILL FILL_2_NAND3X1_17 ( );
FILL FILL_3_NAND3X1_17 ( );
FILL FILL_4_NAND3X1_17 ( );
FILL FILL_5_NAND3X1_17 ( );
FILL FILL_6_NAND3X1_17 ( );
FILL FILL_7_NAND3X1_17 ( );
FILL FILL_8_NAND3X1_17 ( );
FILL FILL_0_NAND3X1_20 ( );
FILL FILL_1_NAND3X1_20 ( );
FILL FILL_2_NAND3X1_20 ( );
FILL FILL_3_NAND3X1_20 ( );
FILL FILL_4_NAND3X1_20 ( );
FILL FILL_5_NAND3X1_20 ( );
FILL FILL_6_NAND3X1_20 ( );
FILL FILL_7_NAND3X1_20 ( );
FILL FILL_8_NAND3X1_20 ( );
FILL FILL_9_NAND3X1_20 ( );
FILL FILL_0_NAND3X1_2 ( );
FILL FILL_1_NAND3X1_2 ( );
FILL FILL_2_NAND3X1_2 ( );
FILL FILL_3_NAND3X1_2 ( );
FILL FILL_4_NAND3X1_2 ( );
FILL FILL_5_NAND3X1_2 ( );
FILL FILL_6_NAND3X1_2 ( );
FILL FILL_7_NAND3X1_2 ( );
FILL FILL_8_NAND3X1_2 ( );
FILL FILL_0_AND2X2_8 ( );
FILL FILL_1_AND2X2_8 ( );
FILL FILL_2_AND2X2_8 ( );
FILL FILL_3_AND2X2_8 ( );
FILL FILL_4_AND2X2_8 ( );
FILL FILL_5_AND2X2_8 ( );
FILL FILL_6_AND2X2_8 ( );
FILL FILL_7_AND2X2_8 ( );
FILL FILL_8_AND2X2_8 ( );
FILL FILL_0_INVX1_23 ( );
FILL FILL_1_INVX1_23 ( );
FILL FILL_2_INVX1_23 ( );
FILL FILL_3_INVX1_23 ( );
FILL FILL_4_INVX1_23 ( );
FILL FILL_0_AND2X2_6 ( );
FILL FILL_1_AND2X2_6 ( );
FILL FILL_2_AND2X2_6 ( );
FILL FILL_3_AND2X2_6 ( );
FILL FILL_4_AND2X2_6 ( );
FILL FILL_5_AND2X2_6 ( );
FILL FILL_6_AND2X2_6 ( );
FILL FILL_7_AND2X2_6 ( );
FILL FILL_8_AND2X2_6 ( );
FILL FILL_9_AND2X2_6 ( );
FILL FILL_0_INVX1_16 ( );
FILL FILL_1_INVX1_16 ( );
FILL FILL_2_INVX1_16 ( );
FILL FILL_3_INVX1_16 ( );
FILL FILL_0_DFFSR_126 ( );
FILL FILL_1_DFFSR_126 ( );
FILL FILL_2_DFFSR_126 ( );
FILL FILL_3_DFFSR_126 ( );
FILL FILL_4_DFFSR_126 ( );
FILL FILL_5_DFFSR_126 ( );
FILL FILL_6_DFFSR_126 ( );
FILL FILL_7_DFFSR_126 ( );
FILL FILL_8_DFFSR_126 ( );
FILL FILL_9_DFFSR_126 ( );
FILL FILL_10_DFFSR_126 ( );
FILL FILL_11_DFFSR_126 ( );
FILL FILL_12_DFFSR_126 ( );
FILL FILL_13_DFFSR_126 ( );
FILL FILL_14_DFFSR_126 ( );
FILL FILL_15_DFFSR_126 ( );
FILL FILL_16_DFFSR_126 ( );
FILL FILL_17_DFFSR_126 ( );
FILL FILL_18_DFFSR_126 ( );
FILL FILL_19_DFFSR_126 ( );
FILL FILL_20_DFFSR_126 ( );
FILL FILL_21_DFFSR_126 ( );
FILL FILL_22_DFFSR_126 ( );
FILL FILL_23_DFFSR_126 ( );
FILL FILL_24_DFFSR_126 ( );
FILL FILL_25_DFFSR_126 ( );
FILL FILL_26_DFFSR_126 ( );
FILL FILL_27_DFFSR_126 ( );
FILL FILL_28_DFFSR_126 ( );
FILL FILL_29_DFFSR_126 ( );
FILL FILL_30_DFFSR_126 ( );
FILL FILL_31_DFFSR_126 ( );
FILL FILL_32_DFFSR_126 ( );
FILL FILL_33_DFFSR_126 ( );
FILL FILL_34_DFFSR_126 ( );
FILL FILL_35_DFFSR_126 ( );
FILL FILL_36_DFFSR_126 ( );
FILL FILL_37_DFFSR_126 ( );
FILL FILL_38_DFFSR_126 ( );
FILL FILL_39_DFFSR_126 ( );
FILL FILL_40_DFFSR_126 ( );
FILL FILL_41_DFFSR_126 ( );
FILL FILL_42_DFFSR_126 ( );
FILL FILL_43_DFFSR_126 ( );
FILL FILL_44_DFFSR_126 ( );
FILL FILL_45_DFFSR_126 ( );
FILL FILL_46_DFFSR_126 ( );
FILL FILL_47_DFFSR_126 ( );
FILL FILL_48_DFFSR_126 ( );
FILL FILL_49_DFFSR_126 ( );
FILL FILL_50_DFFSR_126 ( );
FILL FILL_51_DFFSR_126 ( );
FILL FILL_0_INVX1_9 ( );
FILL FILL_1_INVX1_9 ( );
FILL FILL_2_INVX1_9 ( );
FILL FILL_3_INVX1_9 ( );
FILL FILL_4_INVX1_9 ( );
FILL FILL_0_NAND3X1_123 ( );
FILL FILL_1_NAND3X1_123 ( );
FILL FILL_2_NAND3X1_123 ( );
FILL FILL_3_NAND3X1_123 ( );
FILL FILL_4_NAND3X1_123 ( );
FILL FILL_5_NAND3X1_123 ( );
FILL FILL_6_NAND3X1_123 ( );
FILL FILL_7_NAND3X1_123 ( );
FILL FILL_8_NAND3X1_123 ( );
FILL FILL_0_DFFSR_154 ( );
FILL FILL_1_DFFSR_154 ( );
FILL FILL_2_DFFSR_154 ( );
FILL FILL_3_DFFSR_154 ( );
FILL FILL_4_DFFSR_154 ( );
FILL FILL_5_DFFSR_154 ( );
FILL FILL_6_DFFSR_154 ( );
FILL FILL_7_DFFSR_154 ( );
FILL FILL_8_DFFSR_154 ( );
FILL FILL_9_DFFSR_154 ( );
FILL FILL_10_DFFSR_154 ( );
FILL FILL_11_DFFSR_154 ( );
FILL FILL_12_DFFSR_154 ( );
FILL FILL_13_DFFSR_154 ( );
FILL FILL_14_DFFSR_154 ( );
FILL FILL_15_DFFSR_154 ( );
FILL FILL_16_DFFSR_154 ( );
FILL FILL_17_DFFSR_154 ( );
FILL FILL_18_DFFSR_154 ( );
FILL FILL_19_DFFSR_154 ( );
FILL FILL_20_DFFSR_154 ( );
FILL FILL_21_DFFSR_154 ( );
FILL FILL_22_DFFSR_154 ( );
FILL FILL_23_DFFSR_154 ( );
FILL FILL_24_DFFSR_154 ( );
FILL FILL_25_DFFSR_154 ( );
FILL FILL_26_DFFSR_154 ( );
FILL FILL_27_DFFSR_154 ( );
FILL FILL_28_DFFSR_154 ( );
FILL FILL_29_DFFSR_154 ( );
FILL FILL_30_DFFSR_154 ( );
FILL FILL_31_DFFSR_154 ( );
FILL FILL_32_DFFSR_154 ( );
FILL FILL_33_DFFSR_154 ( );
FILL FILL_34_DFFSR_154 ( );
FILL FILL_35_DFFSR_154 ( );
FILL FILL_36_DFFSR_154 ( );
FILL FILL_37_DFFSR_154 ( );
FILL FILL_38_DFFSR_154 ( );
FILL FILL_39_DFFSR_154 ( );
FILL FILL_40_DFFSR_154 ( );
FILL FILL_41_DFFSR_154 ( );
FILL FILL_42_DFFSR_154 ( );
FILL FILL_43_DFFSR_154 ( );
FILL FILL_44_DFFSR_154 ( );
FILL FILL_45_DFFSR_154 ( );
FILL FILL_46_DFFSR_154 ( );
FILL FILL_47_DFFSR_154 ( );
FILL FILL_48_DFFSR_154 ( );
FILL FILL_49_DFFSR_154 ( );
FILL FILL_50_DFFSR_154 ( );
FILL FILL_0_DFFSR_247 ( );
FILL FILL_1_DFFSR_247 ( );
FILL FILL_2_DFFSR_247 ( );
FILL FILL_3_DFFSR_247 ( );
FILL FILL_4_DFFSR_247 ( );
FILL FILL_5_DFFSR_247 ( );
FILL FILL_6_DFFSR_247 ( );
FILL FILL_7_DFFSR_247 ( );
FILL FILL_8_DFFSR_247 ( );
FILL FILL_9_DFFSR_247 ( );
FILL FILL_10_DFFSR_247 ( );
FILL FILL_11_DFFSR_247 ( );
FILL FILL_12_DFFSR_247 ( );
FILL FILL_13_DFFSR_247 ( );
FILL FILL_14_DFFSR_247 ( );
FILL FILL_15_DFFSR_247 ( );
FILL FILL_16_DFFSR_247 ( );
FILL FILL_17_DFFSR_247 ( );
FILL FILL_18_DFFSR_247 ( );
FILL FILL_19_DFFSR_247 ( );
FILL FILL_20_DFFSR_247 ( );
FILL FILL_21_DFFSR_247 ( );
FILL FILL_22_DFFSR_247 ( );
FILL FILL_23_DFFSR_247 ( );
FILL FILL_24_DFFSR_247 ( );
FILL FILL_25_DFFSR_247 ( );
FILL FILL_26_DFFSR_247 ( );
FILL FILL_27_DFFSR_247 ( );
FILL FILL_28_DFFSR_247 ( );
FILL FILL_29_DFFSR_247 ( );
FILL FILL_30_DFFSR_247 ( );
FILL FILL_31_DFFSR_247 ( );
FILL FILL_32_DFFSR_247 ( );
FILL FILL_33_DFFSR_247 ( );
FILL FILL_34_DFFSR_247 ( );
FILL FILL_35_DFFSR_247 ( );
FILL FILL_36_DFFSR_247 ( );
FILL FILL_37_DFFSR_247 ( );
FILL FILL_38_DFFSR_247 ( );
FILL FILL_39_DFFSR_247 ( );
FILL FILL_40_DFFSR_247 ( );
FILL FILL_41_DFFSR_247 ( );
FILL FILL_42_DFFSR_247 ( );
FILL FILL_43_DFFSR_247 ( );
FILL FILL_44_DFFSR_247 ( );
FILL FILL_45_DFFSR_247 ( );
FILL FILL_46_DFFSR_247 ( );
FILL FILL_47_DFFSR_247 ( );
FILL FILL_48_DFFSR_247 ( );
FILL FILL_49_DFFSR_247 ( );
FILL FILL_50_DFFSR_247 ( );
FILL FILL_0_BUFX2_98 ( );
FILL FILL_1_BUFX2_98 ( );
FILL FILL_2_BUFX2_98 ( );
FILL FILL_3_BUFX2_98 ( );
FILL FILL_4_BUFX2_98 ( );
FILL FILL_5_BUFX2_98 ( );
FILL FILL_6_BUFX2_98 ( );
FILL FILL_0_BUFX2_79 ( );
FILL FILL_1_BUFX2_79 ( );
FILL FILL_2_BUFX2_79 ( );
FILL FILL_3_BUFX2_79 ( );
FILL FILL_4_BUFX2_79 ( );
FILL FILL_5_BUFX2_79 ( );
FILL FILL_6_BUFX2_79 ( );
FILL FILL_0_BUFX2_81 ( );
FILL FILL_1_BUFX2_81 ( );
FILL FILL_2_BUFX2_81 ( );
FILL FILL_3_BUFX2_81 ( );
FILL FILL_4_BUFX2_81 ( );
FILL FILL_5_BUFX2_81 ( );
FILL FILL_6_BUFX2_81 ( );
FILL FILL_0_DFFSR_2 ( );
FILL FILL_1_DFFSR_2 ( );
FILL FILL_2_DFFSR_2 ( );
FILL FILL_3_DFFSR_2 ( );
FILL FILL_4_DFFSR_2 ( );
FILL FILL_5_DFFSR_2 ( );
FILL FILL_6_DFFSR_2 ( );
FILL FILL_7_DFFSR_2 ( );
FILL FILL_8_DFFSR_2 ( );
FILL FILL_9_DFFSR_2 ( );
FILL FILL_10_DFFSR_2 ( );
FILL FILL_11_DFFSR_2 ( );
FILL FILL_12_DFFSR_2 ( );
FILL FILL_13_DFFSR_2 ( );
FILL FILL_14_DFFSR_2 ( );
FILL FILL_15_DFFSR_2 ( );
FILL FILL_16_DFFSR_2 ( );
FILL FILL_17_DFFSR_2 ( );
FILL FILL_18_DFFSR_2 ( );
FILL FILL_19_DFFSR_2 ( );
FILL FILL_20_DFFSR_2 ( );
FILL FILL_21_DFFSR_2 ( );
FILL FILL_22_DFFSR_2 ( );
FILL FILL_23_DFFSR_2 ( );
FILL FILL_24_DFFSR_2 ( );
FILL FILL_25_DFFSR_2 ( );
FILL FILL_26_DFFSR_2 ( );
FILL FILL_27_DFFSR_2 ( );
FILL FILL_28_DFFSR_2 ( );
FILL FILL_29_DFFSR_2 ( );
FILL FILL_30_DFFSR_2 ( );
FILL FILL_31_DFFSR_2 ( );
FILL FILL_32_DFFSR_2 ( );
FILL FILL_33_DFFSR_2 ( );
FILL FILL_34_DFFSR_2 ( );
FILL FILL_35_DFFSR_2 ( );
FILL FILL_36_DFFSR_2 ( );
FILL FILL_37_DFFSR_2 ( );
FILL FILL_38_DFFSR_2 ( );
FILL FILL_39_DFFSR_2 ( );
FILL FILL_40_DFFSR_2 ( );
FILL FILL_41_DFFSR_2 ( );
FILL FILL_42_DFFSR_2 ( );
FILL FILL_43_DFFSR_2 ( );
FILL FILL_44_DFFSR_2 ( );
FILL FILL_45_DFFSR_2 ( );
FILL FILL_46_DFFSR_2 ( );
FILL FILL_47_DFFSR_2 ( );
FILL FILL_48_DFFSR_2 ( );
FILL FILL_49_DFFSR_2 ( );
FILL FILL_50_DFFSR_2 ( );
FILL FILL_0_NAND2X1_155 ( );
FILL FILL_1_NAND2X1_155 ( );
FILL FILL_2_NAND2X1_155 ( );
FILL FILL_3_NAND2X1_155 ( );
FILL FILL_4_NAND2X1_155 ( );
FILL FILL_5_NAND2X1_155 ( );
FILL FILL_6_NAND2X1_155 ( );
FILL FILL_0_AOI21X1_60 ( );
FILL FILL_1_AOI21X1_60 ( );
FILL FILL_2_AOI21X1_60 ( );
FILL FILL_3_AOI21X1_60 ( );
FILL FILL_4_AOI21X1_60 ( );
FILL FILL_5_AOI21X1_60 ( );
FILL FILL_6_AOI21X1_60 ( );
FILL FILL_7_AOI21X1_60 ( );
FILL FILL_8_AOI21X1_60 ( );
FILL FILL_0_CLKBUF1_45 ( );
FILL FILL_1_CLKBUF1_45 ( );
FILL FILL_2_CLKBUF1_45 ( );
FILL FILL_3_CLKBUF1_45 ( );
FILL FILL_4_CLKBUF1_45 ( );
FILL FILL_5_CLKBUF1_45 ( );
FILL FILL_6_CLKBUF1_45 ( );
FILL FILL_7_CLKBUF1_45 ( );
FILL FILL_8_CLKBUF1_45 ( );
FILL FILL_9_CLKBUF1_45 ( );
FILL FILL_10_CLKBUF1_45 ( );
FILL FILL_11_CLKBUF1_45 ( );
FILL FILL_12_CLKBUF1_45 ( );
FILL FILL_13_CLKBUF1_45 ( );
FILL FILL_14_CLKBUF1_45 ( );
FILL FILL_15_CLKBUF1_45 ( );
FILL FILL_16_CLKBUF1_45 ( );
FILL FILL_17_CLKBUF1_45 ( );
FILL FILL_18_CLKBUF1_45 ( );
FILL FILL_19_CLKBUF1_45 ( );
FILL FILL_20_CLKBUF1_45 ( );
FILL FILL_0_DFFSR_76 ( );
FILL FILL_1_DFFSR_76 ( );
FILL FILL_2_DFFSR_76 ( );
FILL FILL_3_DFFSR_76 ( );
FILL FILL_4_DFFSR_76 ( );
FILL FILL_5_DFFSR_76 ( );
FILL FILL_6_DFFSR_76 ( );
FILL FILL_7_DFFSR_76 ( );
FILL FILL_8_DFFSR_76 ( );
FILL FILL_9_DFFSR_76 ( );
FILL FILL_10_DFFSR_76 ( );
FILL FILL_11_DFFSR_76 ( );
FILL FILL_12_DFFSR_76 ( );
FILL FILL_13_DFFSR_76 ( );
FILL FILL_14_DFFSR_76 ( );
FILL FILL_15_DFFSR_76 ( );
FILL FILL_16_DFFSR_76 ( );
FILL FILL_17_DFFSR_76 ( );
FILL FILL_18_DFFSR_76 ( );
FILL FILL_19_DFFSR_76 ( );
FILL FILL_20_DFFSR_76 ( );
FILL FILL_21_DFFSR_76 ( );
FILL FILL_22_DFFSR_76 ( );
FILL FILL_23_DFFSR_76 ( );
FILL FILL_24_DFFSR_76 ( );
FILL FILL_25_DFFSR_76 ( );
FILL FILL_26_DFFSR_76 ( );
FILL FILL_27_DFFSR_76 ( );
FILL FILL_28_DFFSR_76 ( );
FILL FILL_29_DFFSR_76 ( );
FILL FILL_30_DFFSR_76 ( );
FILL FILL_31_DFFSR_76 ( );
FILL FILL_32_DFFSR_76 ( );
FILL FILL_33_DFFSR_76 ( );
FILL FILL_34_DFFSR_76 ( );
FILL FILL_35_DFFSR_76 ( );
FILL FILL_36_DFFSR_76 ( );
FILL FILL_37_DFFSR_76 ( );
FILL FILL_38_DFFSR_76 ( );
FILL FILL_39_DFFSR_76 ( );
FILL FILL_40_DFFSR_76 ( );
FILL FILL_41_DFFSR_76 ( );
FILL FILL_42_DFFSR_76 ( );
FILL FILL_43_DFFSR_76 ( );
FILL FILL_44_DFFSR_76 ( );
FILL FILL_45_DFFSR_76 ( );
FILL FILL_46_DFFSR_76 ( );
FILL FILL_47_DFFSR_76 ( );
FILL FILL_48_DFFSR_76 ( );
FILL FILL_49_DFFSR_76 ( );
FILL FILL_50_DFFSR_76 ( );
FILL FILL_0_NAND3X1_32 ( );
FILL FILL_1_NAND3X1_32 ( );
FILL FILL_2_NAND3X1_32 ( );
FILL FILL_3_NAND3X1_32 ( );
FILL FILL_4_NAND3X1_32 ( );
FILL FILL_5_NAND3X1_32 ( );
FILL FILL_6_NAND3X1_32 ( );
FILL FILL_7_NAND3X1_32 ( );
FILL FILL_8_NAND3X1_32 ( );
FILL FILL_0_NOR2X1_16 ( );
FILL FILL_1_NOR2X1_16 ( );
FILL FILL_2_NOR2X1_16 ( );
FILL FILL_3_NOR2X1_16 ( );
FILL FILL_4_NOR2X1_16 ( );
FILL FILL_5_NOR2X1_16 ( );
FILL FILL_6_NOR2X1_16 ( );
FILL FILL_0_NAND2X1_10 ( );
FILL FILL_1_NAND2X1_10 ( );
FILL FILL_2_NAND2X1_10 ( );
FILL FILL_3_NAND2X1_10 ( );
FILL FILL_4_NAND2X1_10 ( );
FILL FILL_5_NAND2X1_10 ( );
FILL FILL_6_NAND2X1_10 ( );
FILL FILL_0_DFFSR_7 ( );
FILL FILL_1_DFFSR_7 ( );
FILL FILL_2_DFFSR_7 ( );
FILL FILL_3_DFFSR_7 ( );
FILL FILL_4_DFFSR_7 ( );
FILL FILL_5_DFFSR_7 ( );
FILL FILL_6_DFFSR_7 ( );
FILL FILL_7_DFFSR_7 ( );
FILL FILL_8_DFFSR_7 ( );
FILL FILL_9_DFFSR_7 ( );
FILL FILL_10_DFFSR_7 ( );
FILL FILL_11_DFFSR_7 ( );
FILL FILL_12_DFFSR_7 ( );
FILL FILL_13_DFFSR_7 ( );
FILL FILL_14_DFFSR_7 ( );
FILL FILL_15_DFFSR_7 ( );
FILL FILL_16_DFFSR_7 ( );
FILL FILL_17_DFFSR_7 ( );
FILL FILL_18_DFFSR_7 ( );
FILL FILL_19_DFFSR_7 ( );
FILL FILL_20_DFFSR_7 ( );
FILL FILL_21_DFFSR_7 ( );
FILL FILL_22_DFFSR_7 ( );
FILL FILL_23_DFFSR_7 ( );
FILL FILL_24_DFFSR_7 ( );
FILL FILL_25_DFFSR_7 ( );
FILL FILL_26_DFFSR_7 ( );
FILL FILL_27_DFFSR_7 ( );
FILL FILL_28_DFFSR_7 ( );
FILL FILL_29_DFFSR_7 ( );
FILL FILL_30_DFFSR_7 ( );
FILL FILL_31_DFFSR_7 ( );
FILL FILL_32_DFFSR_7 ( );
FILL FILL_33_DFFSR_7 ( );
FILL FILL_34_DFFSR_7 ( );
FILL FILL_35_DFFSR_7 ( );
FILL FILL_36_DFFSR_7 ( );
FILL FILL_37_DFFSR_7 ( );
FILL FILL_38_DFFSR_7 ( );
FILL FILL_39_DFFSR_7 ( );
FILL FILL_40_DFFSR_7 ( );
FILL FILL_41_DFFSR_7 ( );
FILL FILL_42_DFFSR_7 ( );
FILL FILL_43_DFFSR_7 ( );
FILL FILL_44_DFFSR_7 ( );
FILL FILL_45_DFFSR_7 ( );
FILL FILL_46_DFFSR_7 ( );
FILL FILL_47_DFFSR_7 ( );
FILL FILL_48_DFFSR_7 ( );
FILL FILL_49_DFFSR_7 ( );
FILL FILL_50_DFFSR_7 ( );
FILL FILL_0_DFFSR_65 ( );
FILL FILL_1_DFFSR_65 ( );
FILL FILL_2_DFFSR_65 ( );
FILL FILL_3_DFFSR_65 ( );
FILL FILL_4_DFFSR_65 ( );
FILL FILL_5_DFFSR_65 ( );
FILL FILL_6_DFFSR_65 ( );
FILL FILL_7_DFFSR_65 ( );
FILL FILL_8_DFFSR_65 ( );
FILL FILL_9_DFFSR_65 ( );
FILL FILL_10_DFFSR_65 ( );
FILL FILL_11_DFFSR_65 ( );
FILL FILL_12_DFFSR_65 ( );
FILL FILL_13_DFFSR_65 ( );
FILL FILL_14_DFFSR_65 ( );
FILL FILL_15_DFFSR_65 ( );
FILL FILL_16_DFFSR_65 ( );
FILL FILL_17_DFFSR_65 ( );
FILL FILL_18_DFFSR_65 ( );
FILL FILL_19_DFFSR_65 ( );
FILL FILL_20_DFFSR_65 ( );
FILL FILL_21_DFFSR_65 ( );
FILL FILL_22_DFFSR_65 ( );
FILL FILL_23_DFFSR_65 ( );
FILL FILL_24_DFFSR_65 ( );
FILL FILL_25_DFFSR_65 ( );
FILL FILL_26_DFFSR_65 ( );
FILL FILL_27_DFFSR_65 ( );
FILL FILL_28_DFFSR_65 ( );
FILL FILL_29_DFFSR_65 ( );
FILL FILL_30_DFFSR_65 ( );
FILL FILL_31_DFFSR_65 ( );
FILL FILL_32_DFFSR_65 ( );
FILL FILL_33_DFFSR_65 ( );
FILL FILL_34_DFFSR_65 ( );
FILL FILL_35_DFFSR_65 ( );
FILL FILL_36_DFFSR_65 ( );
FILL FILL_37_DFFSR_65 ( );
FILL FILL_38_DFFSR_65 ( );
FILL FILL_39_DFFSR_65 ( );
FILL FILL_40_DFFSR_65 ( );
FILL FILL_41_DFFSR_65 ( );
FILL FILL_42_DFFSR_65 ( );
FILL FILL_43_DFFSR_65 ( );
FILL FILL_44_DFFSR_65 ( );
FILL FILL_45_DFFSR_65 ( );
FILL FILL_46_DFFSR_65 ( );
FILL FILL_47_DFFSR_65 ( );
FILL FILL_48_DFFSR_65 ( );
FILL FILL_49_DFFSR_65 ( );
FILL FILL_50_DFFSR_65 ( );
FILL FILL_0_NAND2X1_16 ( );
FILL FILL_1_NAND2X1_16 ( );
FILL FILL_2_NAND2X1_16 ( );
FILL FILL_3_NAND2X1_16 ( );
FILL FILL_4_NAND2X1_16 ( );
FILL FILL_5_NAND2X1_16 ( );
FILL FILL_6_NAND2X1_16 ( );
FILL FILL_0_NAND3X1_18 ( );
FILL FILL_1_NAND3X1_18 ( );
FILL FILL_2_NAND3X1_18 ( );
FILL FILL_3_NAND3X1_18 ( );
FILL FILL_4_NAND3X1_18 ( );
FILL FILL_5_NAND3X1_18 ( );
FILL FILL_6_NAND3X1_18 ( );
FILL FILL_7_NAND3X1_18 ( );
FILL FILL_8_NAND3X1_18 ( );
FILL FILL_9_NAND3X1_18 ( );
FILL FILL_0_OAI21X1_2 ( );
FILL FILL_1_OAI21X1_2 ( );
FILL FILL_2_OAI21X1_2 ( );
FILL FILL_3_OAI21X1_2 ( );
FILL FILL_4_OAI21X1_2 ( );
FILL FILL_5_OAI21X1_2 ( );
FILL FILL_6_OAI21X1_2 ( );
FILL FILL_7_OAI21X1_2 ( );
FILL FILL_8_OAI21X1_2 ( );
FILL FILL_9_OAI21X1_2 ( );
FILL FILL_0_OAI21X1_1 ( );
FILL FILL_1_OAI21X1_1 ( );
FILL FILL_2_OAI21X1_1 ( );
FILL FILL_3_OAI21X1_1 ( );
FILL FILL_4_OAI21X1_1 ( );
FILL FILL_5_OAI21X1_1 ( );
FILL FILL_6_OAI21X1_1 ( );
FILL FILL_7_OAI21X1_1 ( );
FILL FILL_8_OAI21X1_1 ( );
FILL FILL_9_OAI21X1_1 ( );
FILL FILL_0_NAND3X1_4 ( );
FILL FILL_1_NAND3X1_4 ( );
FILL FILL_2_NAND3X1_4 ( );
FILL FILL_3_NAND3X1_4 ( );
FILL FILL_4_NAND3X1_4 ( );
FILL FILL_5_NAND3X1_4 ( );
FILL FILL_6_NAND3X1_4 ( );
FILL FILL_7_NAND3X1_4 ( );
FILL FILL_8_NAND3X1_4 ( );
FILL FILL_0_DFFSR_122 ( );
FILL FILL_1_DFFSR_122 ( );
FILL FILL_2_DFFSR_122 ( );
FILL FILL_3_DFFSR_122 ( );
FILL FILL_4_DFFSR_122 ( );
FILL FILL_5_DFFSR_122 ( );
FILL FILL_6_DFFSR_122 ( );
FILL FILL_7_DFFSR_122 ( );
FILL FILL_8_DFFSR_122 ( );
FILL FILL_9_DFFSR_122 ( );
FILL FILL_10_DFFSR_122 ( );
FILL FILL_11_DFFSR_122 ( );
FILL FILL_12_DFFSR_122 ( );
FILL FILL_13_DFFSR_122 ( );
FILL FILL_14_DFFSR_122 ( );
FILL FILL_15_DFFSR_122 ( );
FILL FILL_16_DFFSR_122 ( );
FILL FILL_17_DFFSR_122 ( );
FILL FILL_18_DFFSR_122 ( );
FILL FILL_19_DFFSR_122 ( );
FILL FILL_20_DFFSR_122 ( );
FILL FILL_21_DFFSR_122 ( );
FILL FILL_22_DFFSR_122 ( );
FILL FILL_23_DFFSR_122 ( );
FILL FILL_24_DFFSR_122 ( );
FILL FILL_25_DFFSR_122 ( );
FILL FILL_26_DFFSR_122 ( );
FILL FILL_27_DFFSR_122 ( );
FILL FILL_28_DFFSR_122 ( );
FILL FILL_29_DFFSR_122 ( );
FILL FILL_30_DFFSR_122 ( );
FILL FILL_31_DFFSR_122 ( );
FILL FILL_32_DFFSR_122 ( );
FILL FILL_33_DFFSR_122 ( );
FILL FILL_34_DFFSR_122 ( );
FILL FILL_35_DFFSR_122 ( );
FILL FILL_36_DFFSR_122 ( );
FILL FILL_37_DFFSR_122 ( );
FILL FILL_38_DFFSR_122 ( );
FILL FILL_39_DFFSR_122 ( );
FILL FILL_40_DFFSR_122 ( );
FILL FILL_41_DFFSR_122 ( );
FILL FILL_42_DFFSR_122 ( );
FILL FILL_43_DFFSR_122 ( );
FILL FILL_44_DFFSR_122 ( );
FILL FILL_45_DFFSR_122 ( );
FILL FILL_46_DFFSR_122 ( );
FILL FILL_47_DFFSR_122 ( );
FILL FILL_48_DFFSR_122 ( );
FILL FILL_49_DFFSR_122 ( );
FILL FILL_50_DFFSR_122 ( );
FILL FILL_0_BUFX2_83 ( );
FILL FILL_1_BUFX2_83 ( );
FILL FILL_2_BUFX2_83 ( );
FILL FILL_3_BUFX2_83 ( );
FILL FILL_4_BUFX2_83 ( );
FILL FILL_5_BUFX2_83 ( );
FILL FILL_6_BUFX2_83 ( );
FILL FILL_0_NAND3X1_115 ( );
FILL FILL_1_NAND3X1_115 ( );
FILL FILL_2_NAND3X1_115 ( );
FILL FILL_3_NAND3X1_115 ( );
FILL FILL_4_NAND3X1_115 ( );
FILL FILL_5_NAND3X1_115 ( );
FILL FILL_6_NAND3X1_115 ( );
FILL FILL_7_NAND3X1_115 ( );
FILL FILL_8_NAND3X1_115 ( );
FILL FILL_9_NAND3X1_115 ( );
FILL FILL_0_NAND3X1_75 ( );
FILL FILL_1_NAND3X1_75 ( );
FILL FILL_2_NAND3X1_75 ( );
FILL FILL_3_NAND3X1_75 ( );
FILL FILL_4_NAND3X1_75 ( );
FILL FILL_5_NAND3X1_75 ( );
FILL FILL_6_NAND3X1_75 ( );
FILL FILL_7_NAND3X1_75 ( );
FILL FILL_8_NAND3X1_75 ( );
FILL FILL_0_OAI21X1_10 ( );
FILL FILL_1_OAI21X1_10 ( );
FILL FILL_2_OAI21X1_10 ( );
FILL FILL_3_OAI21X1_10 ( );
FILL FILL_4_OAI21X1_10 ( );
FILL FILL_5_OAI21X1_10 ( );
FILL FILL_6_OAI21X1_10 ( );
FILL FILL_7_OAI21X1_10 ( );
FILL FILL_8_OAI21X1_10 ( );
FILL FILL_0_DFFSR_146 ( );
FILL FILL_1_DFFSR_146 ( );
FILL FILL_2_DFFSR_146 ( );
FILL FILL_3_DFFSR_146 ( );
FILL FILL_4_DFFSR_146 ( );
FILL FILL_5_DFFSR_146 ( );
FILL FILL_6_DFFSR_146 ( );
FILL FILL_7_DFFSR_146 ( );
FILL FILL_8_DFFSR_146 ( );
FILL FILL_9_DFFSR_146 ( );
FILL FILL_10_DFFSR_146 ( );
FILL FILL_11_DFFSR_146 ( );
FILL FILL_12_DFFSR_146 ( );
FILL FILL_13_DFFSR_146 ( );
FILL FILL_14_DFFSR_146 ( );
FILL FILL_15_DFFSR_146 ( );
FILL FILL_16_DFFSR_146 ( );
FILL FILL_17_DFFSR_146 ( );
FILL FILL_18_DFFSR_146 ( );
FILL FILL_19_DFFSR_146 ( );
FILL FILL_20_DFFSR_146 ( );
FILL FILL_21_DFFSR_146 ( );
FILL FILL_22_DFFSR_146 ( );
FILL FILL_23_DFFSR_146 ( );
FILL FILL_24_DFFSR_146 ( );
FILL FILL_25_DFFSR_146 ( );
FILL FILL_26_DFFSR_146 ( );
FILL FILL_27_DFFSR_146 ( );
FILL FILL_28_DFFSR_146 ( );
FILL FILL_29_DFFSR_146 ( );
FILL FILL_30_DFFSR_146 ( );
FILL FILL_31_DFFSR_146 ( );
FILL FILL_32_DFFSR_146 ( );
FILL FILL_33_DFFSR_146 ( );
FILL FILL_34_DFFSR_146 ( );
FILL FILL_35_DFFSR_146 ( );
FILL FILL_36_DFFSR_146 ( );
FILL FILL_37_DFFSR_146 ( );
FILL FILL_38_DFFSR_146 ( );
FILL FILL_39_DFFSR_146 ( );
FILL FILL_40_DFFSR_146 ( );
FILL FILL_41_DFFSR_146 ( );
FILL FILL_42_DFFSR_146 ( );
FILL FILL_43_DFFSR_146 ( );
FILL FILL_44_DFFSR_146 ( );
FILL FILL_45_DFFSR_146 ( );
FILL FILL_46_DFFSR_146 ( );
FILL FILL_47_DFFSR_146 ( );
FILL FILL_48_DFFSR_146 ( );
FILL FILL_49_DFFSR_146 ( );
FILL FILL_50_DFFSR_146 ( );
FILL FILL_51_DFFSR_146 ( );
FILL FILL_0_OAI21X1_87 ( );
FILL FILL_1_OAI21X1_87 ( );
FILL FILL_2_OAI21X1_87 ( );
FILL FILL_3_OAI21X1_87 ( );
FILL FILL_4_OAI21X1_87 ( );
FILL FILL_5_OAI21X1_87 ( );
FILL FILL_6_OAI21X1_87 ( );
FILL FILL_7_OAI21X1_87 ( );
FILL FILL_8_OAI21X1_87 ( );
FILL FILL_0_BUFX2_80 ( );
FILL FILL_1_BUFX2_80 ( );
FILL FILL_2_BUFX2_80 ( );
FILL FILL_3_BUFX2_80 ( );
FILL FILL_4_BUFX2_80 ( );
FILL FILL_5_BUFX2_80 ( );
FILL FILL_6_BUFX2_80 ( );
FILL FILL_0_BUFX2_100 ( );
FILL FILL_1_BUFX2_100 ( );
FILL FILL_2_BUFX2_100 ( );
FILL FILL_3_BUFX2_100 ( );
FILL FILL_4_BUFX2_100 ( );
FILL FILL_5_BUFX2_100 ( );
FILL FILL_6_BUFX2_100 ( );
FILL FILL_0_INVX1_186 ( );
FILL FILL_1_INVX1_186 ( );
FILL FILL_2_INVX1_186 ( );
FILL FILL_3_INVX1_186 ( );
FILL FILL_4_INVX1_186 ( );
FILL FILL_0_DFFSR_6 ( );
FILL FILL_1_DFFSR_6 ( );
FILL FILL_2_DFFSR_6 ( );
FILL FILL_3_DFFSR_6 ( );
FILL FILL_4_DFFSR_6 ( );
FILL FILL_5_DFFSR_6 ( );
FILL FILL_6_DFFSR_6 ( );
FILL FILL_7_DFFSR_6 ( );
FILL FILL_8_DFFSR_6 ( );
FILL FILL_9_DFFSR_6 ( );
FILL FILL_10_DFFSR_6 ( );
FILL FILL_11_DFFSR_6 ( );
FILL FILL_12_DFFSR_6 ( );
FILL FILL_13_DFFSR_6 ( );
FILL FILL_14_DFFSR_6 ( );
FILL FILL_15_DFFSR_6 ( );
FILL FILL_16_DFFSR_6 ( );
FILL FILL_17_DFFSR_6 ( );
FILL FILL_18_DFFSR_6 ( );
FILL FILL_19_DFFSR_6 ( );
FILL FILL_20_DFFSR_6 ( );
FILL FILL_21_DFFSR_6 ( );
FILL FILL_22_DFFSR_6 ( );
FILL FILL_23_DFFSR_6 ( );
FILL FILL_24_DFFSR_6 ( );
FILL FILL_25_DFFSR_6 ( );
FILL FILL_26_DFFSR_6 ( );
FILL FILL_27_DFFSR_6 ( );
FILL FILL_28_DFFSR_6 ( );
FILL FILL_29_DFFSR_6 ( );
FILL FILL_30_DFFSR_6 ( );
FILL FILL_31_DFFSR_6 ( );
FILL FILL_32_DFFSR_6 ( );
FILL FILL_33_DFFSR_6 ( );
FILL FILL_34_DFFSR_6 ( );
FILL FILL_35_DFFSR_6 ( );
FILL FILL_36_DFFSR_6 ( );
FILL FILL_37_DFFSR_6 ( );
FILL FILL_38_DFFSR_6 ( );
FILL FILL_39_DFFSR_6 ( );
FILL FILL_40_DFFSR_6 ( );
FILL FILL_41_DFFSR_6 ( );
FILL FILL_42_DFFSR_6 ( );
FILL FILL_43_DFFSR_6 ( );
FILL FILL_44_DFFSR_6 ( );
FILL FILL_45_DFFSR_6 ( );
FILL FILL_46_DFFSR_6 ( );
FILL FILL_47_DFFSR_6 ( );
FILL FILL_48_DFFSR_6 ( );
FILL FILL_49_DFFSR_6 ( );
FILL FILL_50_DFFSR_6 ( );
FILL FILL_51_DFFSR_6 ( );
FILL FILL_0_DFFPOSX1_25 ( );
FILL FILL_1_DFFPOSX1_25 ( );
FILL FILL_2_DFFPOSX1_25 ( );
FILL FILL_3_DFFPOSX1_25 ( );
FILL FILL_4_DFFPOSX1_25 ( );
FILL FILL_5_DFFPOSX1_25 ( );
FILL FILL_6_DFFPOSX1_25 ( );
FILL FILL_7_DFFPOSX1_25 ( );
FILL FILL_8_DFFPOSX1_25 ( );
FILL FILL_9_DFFPOSX1_25 ( );
FILL FILL_10_DFFPOSX1_25 ( );
FILL FILL_11_DFFPOSX1_25 ( );
FILL FILL_12_DFFPOSX1_25 ( );
FILL FILL_13_DFFPOSX1_25 ( );
FILL FILL_14_DFFPOSX1_25 ( );
FILL FILL_15_DFFPOSX1_25 ( );
FILL FILL_16_DFFPOSX1_25 ( );
FILL FILL_17_DFFPOSX1_25 ( );
FILL FILL_18_DFFPOSX1_25 ( );
FILL FILL_19_DFFPOSX1_25 ( );
FILL FILL_20_DFFPOSX1_25 ( );
FILL FILL_21_DFFPOSX1_25 ( );
FILL FILL_22_DFFPOSX1_25 ( );
FILL FILL_23_DFFPOSX1_25 ( );
FILL FILL_24_DFFPOSX1_25 ( );
FILL FILL_25_DFFPOSX1_25 ( );
FILL FILL_26_DFFPOSX1_25 ( );
FILL FILL_27_DFFPOSX1_25 ( );
FILL FILL_0_NAND2X1_168 ( );
FILL FILL_1_NAND2X1_168 ( );
FILL FILL_2_NAND2X1_168 ( );
FILL FILL_3_NAND2X1_168 ( );
FILL FILL_4_NAND2X1_168 ( );
FILL FILL_5_NAND2X1_168 ( );
FILL FILL_6_NAND2X1_168 ( );
FILL FILL_0_DFFSR_26 ( );
FILL FILL_1_DFFSR_26 ( );
FILL FILL_2_DFFSR_26 ( );
FILL FILL_3_DFFSR_26 ( );
FILL FILL_4_DFFSR_26 ( );
FILL FILL_5_DFFSR_26 ( );
FILL FILL_6_DFFSR_26 ( );
FILL FILL_7_DFFSR_26 ( );
FILL FILL_8_DFFSR_26 ( );
FILL FILL_9_DFFSR_26 ( );
FILL FILL_10_DFFSR_26 ( );
FILL FILL_11_DFFSR_26 ( );
FILL FILL_12_DFFSR_26 ( );
FILL FILL_13_DFFSR_26 ( );
FILL FILL_14_DFFSR_26 ( );
FILL FILL_15_DFFSR_26 ( );
FILL FILL_16_DFFSR_26 ( );
FILL FILL_17_DFFSR_26 ( );
FILL FILL_18_DFFSR_26 ( );
FILL FILL_19_DFFSR_26 ( );
FILL FILL_20_DFFSR_26 ( );
FILL FILL_21_DFFSR_26 ( );
FILL FILL_22_DFFSR_26 ( );
FILL FILL_23_DFFSR_26 ( );
FILL FILL_24_DFFSR_26 ( );
FILL FILL_25_DFFSR_26 ( );
FILL FILL_26_DFFSR_26 ( );
FILL FILL_27_DFFSR_26 ( );
FILL FILL_28_DFFSR_26 ( );
FILL FILL_29_DFFSR_26 ( );
FILL FILL_30_DFFSR_26 ( );
FILL FILL_31_DFFSR_26 ( );
FILL FILL_32_DFFSR_26 ( );
FILL FILL_33_DFFSR_26 ( );
FILL FILL_34_DFFSR_26 ( );
FILL FILL_35_DFFSR_26 ( );
FILL FILL_36_DFFSR_26 ( );
FILL FILL_37_DFFSR_26 ( );
FILL FILL_38_DFFSR_26 ( );
FILL FILL_39_DFFSR_26 ( );
FILL FILL_40_DFFSR_26 ( );
FILL FILL_41_DFFSR_26 ( );
FILL FILL_42_DFFSR_26 ( );
FILL FILL_43_DFFSR_26 ( );
FILL FILL_44_DFFSR_26 ( );
FILL FILL_45_DFFSR_26 ( );
FILL FILL_46_DFFSR_26 ( );
FILL FILL_47_DFFSR_26 ( );
FILL FILL_48_DFFSR_26 ( );
FILL FILL_49_DFFSR_26 ( );
FILL FILL_50_DFFSR_26 ( );
FILL FILL_0_NOR2X1_17 ( );
FILL FILL_1_NOR2X1_17 ( );
FILL FILL_2_NOR2X1_17 ( );
FILL FILL_3_NOR2X1_17 ( );
FILL FILL_4_NOR2X1_17 ( );
FILL FILL_5_NOR2X1_17 ( );
FILL FILL_6_NOR2X1_17 ( );
FILL FILL_0_NAND3X1_31 ( );
FILL FILL_1_NAND3X1_31 ( );
FILL FILL_2_NAND3X1_31 ( );
FILL FILL_3_NAND3X1_31 ( );
FILL FILL_4_NAND3X1_31 ( );
FILL FILL_5_NAND3X1_31 ( );
FILL FILL_6_NAND3X1_31 ( );
FILL FILL_7_NAND3X1_31 ( );
FILL FILL_8_NAND3X1_31 ( );
FILL FILL_0_NAND3X1_30 ( );
FILL FILL_1_NAND3X1_30 ( );
FILL FILL_2_NAND3X1_30 ( );
FILL FILL_3_NAND3X1_30 ( );
FILL FILL_4_NAND3X1_30 ( );
FILL FILL_5_NAND3X1_30 ( );
FILL FILL_6_NAND3X1_30 ( );
FILL FILL_7_NAND3X1_30 ( );
FILL FILL_8_NAND3X1_30 ( );
FILL FILL_0_NAND3X1_42 ( );
FILL FILL_1_NAND3X1_42 ( );
FILL FILL_2_NAND3X1_42 ( );
FILL FILL_3_NAND3X1_42 ( );
FILL FILL_4_NAND3X1_42 ( );
FILL FILL_5_NAND3X1_42 ( );
FILL FILL_6_NAND3X1_42 ( );
FILL FILL_7_NAND3X1_42 ( );
FILL FILL_8_NAND3X1_42 ( );
FILL FILL_9_NAND3X1_42 ( );
FILL FILL_0_NAND3X1_10 ( );
FILL FILL_1_NAND3X1_10 ( );
FILL FILL_2_NAND3X1_10 ( );
FILL FILL_3_NAND3X1_10 ( );
FILL FILL_4_NAND3X1_10 ( );
FILL FILL_5_NAND3X1_10 ( );
FILL FILL_6_NAND3X1_10 ( );
FILL FILL_7_NAND3X1_10 ( );
FILL FILL_8_NAND3X1_10 ( );
FILL FILL_0_DFFSR_31 ( );
FILL FILL_1_DFFSR_31 ( );
FILL FILL_2_DFFSR_31 ( );
FILL FILL_3_DFFSR_31 ( );
FILL FILL_4_DFFSR_31 ( );
FILL FILL_5_DFFSR_31 ( );
FILL FILL_6_DFFSR_31 ( );
FILL FILL_7_DFFSR_31 ( );
FILL FILL_8_DFFSR_31 ( );
FILL FILL_9_DFFSR_31 ( );
FILL FILL_10_DFFSR_31 ( );
FILL FILL_11_DFFSR_31 ( );
FILL FILL_12_DFFSR_31 ( );
FILL FILL_13_DFFSR_31 ( );
FILL FILL_14_DFFSR_31 ( );
FILL FILL_15_DFFSR_31 ( );
FILL FILL_16_DFFSR_31 ( );
FILL FILL_17_DFFSR_31 ( );
FILL FILL_18_DFFSR_31 ( );
FILL FILL_19_DFFSR_31 ( );
FILL FILL_20_DFFSR_31 ( );
FILL FILL_21_DFFSR_31 ( );
FILL FILL_22_DFFSR_31 ( );
FILL FILL_23_DFFSR_31 ( );
FILL FILL_24_DFFSR_31 ( );
FILL FILL_25_DFFSR_31 ( );
FILL FILL_26_DFFSR_31 ( );
FILL FILL_27_DFFSR_31 ( );
FILL FILL_28_DFFSR_31 ( );
FILL FILL_29_DFFSR_31 ( );
FILL FILL_30_DFFSR_31 ( );
FILL FILL_31_DFFSR_31 ( );
FILL FILL_32_DFFSR_31 ( );
FILL FILL_33_DFFSR_31 ( );
FILL FILL_34_DFFSR_31 ( );
FILL FILL_35_DFFSR_31 ( );
FILL FILL_36_DFFSR_31 ( );
FILL FILL_37_DFFSR_31 ( );
FILL FILL_38_DFFSR_31 ( );
FILL FILL_39_DFFSR_31 ( );
FILL FILL_40_DFFSR_31 ( );
FILL FILL_41_DFFSR_31 ( );
FILL FILL_42_DFFSR_31 ( );
FILL FILL_43_DFFSR_31 ( );
FILL FILL_44_DFFSR_31 ( );
FILL FILL_45_DFFSR_31 ( );
FILL FILL_46_DFFSR_31 ( );
FILL FILL_47_DFFSR_31 ( );
FILL FILL_48_DFFSR_31 ( );
FILL FILL_49_DFFSR_31 ( );
FILL FILL_50_DFFSR_31 ( );
FILL FILL_0_DFFSR_9 ( );
FILL FILL_1_DFFSR_9 ( );
FILL FILL_2_DFFSR_9 ( );
FILL FILL_3_DFFSR_9 ( );
FILL FILL_4_DFFSR_9 ( );
FILL FILL_5_DFFSR_9 ( );
FILL FILL_6_DFFSR_9 ( );
FILL FILL_7_DFFSR_9 ( );
FILL FILL_8_DFFSR_9 ( );
FILL FILL_9_DFFSR_9 ( );
FILL FILL_10_DFFSR_9 ( );
FILL FILL_11_DFFSR_9 ( );
FILL FILL_12_DFFSR_9 ( );
FILL FILL_13_DFFSR_9 ( );
FILL FILL_14_DFFSR_9 ( );
FILL FILL_15_DFFSR_9 ( );
FILL FILL_16_DFFSR_9 ( );
FILL FILL_17_DFFSR_9 ( );
FILL FILL_18_DFFSR_9 ( );
FILL FILL_19_DFFSR_9 ( );
FILL FILL_20_DFFSR_9 ( );
FILL FILL_21_DFFSR_9 ( );
FILL FILL_22_DFFSR_9 ( );
FILL FILL_23_DFFSR_9 ( );
FILL FILL_24_DFFSR_9 ( );
FILL FILL_25_DFFSR_9 ( );
FILL FILL_26_DFFSR_9 ( );
FILL FILL_27_DFFSR_9 ( );
FILL FILL_28_DFFSR_9 ( );
FILL FILL_29_DFFSR_9 ( );
FILL FILL_30_DFFSR_9 ( );
FILL FILL_31_DFFSR_9 ( );
FILL FILL_32_DFFSR_9 ( );
FILL FILL_33_DFFSR_9 ( );
FILL FILL_34_DFFSR_9 ( );
FILL FILL_35_DFFSR_9 ( );
FILL FILL_36_DFFSR_9 ( );
FILL FILL_37_DFFSR_9 ( );
FILL FILL_38_DFFSR_9 ( );
FILL FILL_39_DFFSR_9 ( );
FILL FILL_40_DFFSR_9 ( );
FILL FILL_41_DFFSR_9 ( );
FILL FILL_42_DFFSR_9 ( );
FILL FILL_43_DFFSR_9 ( );
FILL FILL_44_DFFSR_9 ( );
FILL FILL_45_DFFSR_9 ( );
FILL FILL_46_DFFSR_9 ( );
FILL FILL_47_DFFSR_9 ( );
FILL FILL_48_DFFSR_9 ( );
FILL FILL_49_DFFSR_9 ( );
FILL FILL_50_DFFSR_9 ( );
FILL FILL_0_NAND2X1_9 ( );
FILL FILL_1_NAND2X1_9 ( );
FILL FILL_2_NAND2X1_9 ( );
FILL FILL_3_NAND2X1_9 ( );
FILL FILL_4_NAND2X1_9 ( );
FILL FILL_5_NAND2X1_9 ( );
FILL FILL_6_NAND2X1_9 ( );
FILL FILL_0_DFFSR_57 ( );
FILL FILL_1_DFFSR_57 ( );
FILL FILL_2_DFFSR_57 ( );
FILL FILL_3_DFFSR_57 ( );
FILL FILL_4_DFFSR_57 ( );
FILL FILL_5_DFFSR_57 ( );
FILL FILL_6_DFFSR_57 ( );
FILL FILL_7_DFFSR_57 ( );
FILL FILL_8_DFFSR_57 ( );
FILL FILL_9_DFFSR_57 ( );
FILL FILL_10_DFFSR_57 ( );
FILL FILL_11_DFFSR_57 ( );
FILL FILL_12_DFFSR_57 ( );
FILL FILL_13_DFFSR_57 ( );
FILL FILL_14_DFFSR_57 ( );
FILL FILL_15_DFFSR_57 ( );
FILL FILL_16_DFFSR_57 ( );
FILL FILL_17_DFFSR_57 ( );
FILL FILL_18_DFFSR_57 ( );
FILL FILL_19_DFFSR_57 ( );
FILL FILL_20_DFFSR_57 ( );
FILL FILL_21_DFFSR_57 ( );
FILL FILL_22_DFFSR_57 ( );
FILL FILL_23_DFFSR_57 ( );
FILL FILL_24_DFFSR_57 ( );
FILL FILL_25_DFFSR_57 ( );
FILL FILL_26_DFFSR_57 ( );
FILL FILL_27_DFFSR_57 ( );
FILL FILL_28_DFFSR_57 ( );
FILL FILL_29_DFFSR_57 ( );
FILL FILL_30_DFFSR_57 ( );
FILL FILL_31_DFFSR_57 ( );
FILL FILL_32_DFFSR_57 ( );
FILL FILL_33_DFFSR_57 ( );
FILL FILL_34_DFFSR_57 ( );
FILL FILL_35_DFFSR_57 ( );
FILL FILL_36_DFFSR_57 ( );
FILL FILL_37_DFFSR_57 ( );
FILL FILL_38_DFFSR_57 ( );
FILL FILL_39_DFFSR_57 ( );
FILL FILL_40_DFFSR_57 ( );
FILL FILL_41_DFFSR_57 ( );
FILL FILL_42_DFFSR_57 ( );
FILL FILL_43_DFFSR_57 ( );
FILL FILL_44_DFFSR_57 ( );
FILL FILL_45_DFFSR_57 ( );
FILL FILL_46_DFFSR_57 ( );
FILL FILL_47_DFFSR_57 ( );
FILL FILL_48_DFFSR_57 ( );
FILL FILL_49_DFFSR_57 ( );
FILL FILL_50_DFFSR_57 ( );
FILL FILL_51_DFFSR_57 ( );
FILL FILL_0_BUFX2_6 ( );
FILL FILL_1_BUFX2_6 ( );
FILL FILL_2_BUFX2_6 ( );
FILL FILL_3_BUFX2_6 ( );
FILL FILL_4_BUFX2_6 ( );
FILL FILL_5_BUFX2_6 ( );
FILL FILL_6_BUFX2_6 ( );
FILL FILL_0_DFFSR_130 ( );
FILL FILL_1_DFFSR_130 ( );
FILL FILL_2_DFFSR_130 ( );
FILL FILL_3_DFFSR_130 ( );
FILL FILL_4_DFFSR_130 ( );
FILL FILL_5_DFFSR_130 ( );
FILL FILL_6_DFFSR_130 ( );
FILL FILL_7_DFFSR_130 ( );
FILL FILL_8_DFFSR_130 ( );
FILL FILL_9_DFFSR_130 ( );
FILL FILL_10_DFFSR_130 ( );
FILL FILL_11_DFFSR_130 ( );
FILL FILL_12_DFFSR_130 ( );
FILL FILL_13_DFFSR_130 ( );
FILL FILL_14_DFFSR_130 ( );
FILL FILL_15_DFFSR_130 ( );
FILL FILL_16_DFFSR_130 ( );
FILL FILL_17_DFFSR_130 ( );
FILL FILL_18_DFFSR_130 ( );
FILL FILL_19_DFFSR_130 ( );
FILL FILL_20_DFFSR_130 ( );
FILL FILL_21_DFFSR_130 ( );
FILL FILL_22_DFFSR_130 ( );
FILL FILL_23_DFFSR_130 ( );
FILL FILL_24_DFFSR_130 ( );
FILL FILL_25_DFFSR_130 ( );
FILL FILL_26_DFFSR_130 ( );
FILL FILL_27_DFFSR_130 ( );
FILL FILL_28_DFFSR_130 ( );
FILL FILL_29_DFFSR_130 ( );
FILL FILL_30_DFFSR_130 ( );
FILL FILL_31_DFFSR_130 ( );
FILL FILL_32_DFFSR_130 ( );
FILL FILL_33_DFFSR_130 ( );
FILL FILL_34_DFFSR_130 ( );
FILL FILL_35_DFFSR_130 ( );
FILL FILL_36_DFFSR_130 ( );
FILL FILL_37_DFFSR_130 ( );
FILL FILL_38_DFFSR_130 ( );
FILL FILL_39_DFFSR_130 ( );
FILL FILL_40_DFFSR_130 ( );
FILL FILL_41_DFFSR_130 ( );
FILL FILL_42_DFFSR_130 ( );
FILL FILL_43_DFFSR_130 ( );
FILL FILL_44_DFFSR_130 ( );
FILL FILL_45_DFFSR_130 ( );
FILL FILL_46_DFFSR_130 ( );
FILL FILL_47_DFFSR_130 ( );
FILL FILL_48_DFFSR_130 ( );
FILL FILL_49_DFFSR_130 ( );
FILL FILL_50_DFFSR_130 ( );
FILL FILL_0_INVX1_71 ( );
FILL FILL_1_INVX1_71 ( );
FILL FILL_2_INVX1_71 ( );
FILL FILL_3_INVX1_71 ( );
FILL FILL_4_INVX1_71 ( );
FILL FILL_0_DFFSR_259 ( );
FILL FILL_1_DFFSR_259 ( );
FILL FILL_2_DFFSR_259 ( );
FILL FILL_3_DFFSR_259 ( );
FILL FILL_4_DFFSR_259 ( );
FILL FILL_5_DFFSR_259 ( );
FILL FILL_6_DFFSR_259 ( );
FILL FILL_7_DFFSR_259 ( );
FILL FILL_8_DFFSR_259 ( );
FILL FILL_9_DFFSR_259 ( );
FILL FILL_10_DFFSR_259 ( );
FILL FILL_11_DFFSR_259 ( );
FILL FILL_12_DFFSR_259 ( );
FILL FILL_13_DFFSR_259 ( );
FILL FILL_14_DFFSR_259 ( );
FILL FILL_15_DFFSR_259 ( );
FILL FILL_16_DFFSR_259 ( );
FILL FILL_17_DFFSR_259 ( );
FILL FILL_18_DFFSR_259 ( );
FILL FILL_19_DFFSR_259 ( );
FILL FILL_20_DFFSR_259 ( );
FILL FILL_21_DFFSR_259 ( );
FILL FILL_22_DFFSR_259 ( );
FILL FILL_23_DFFSR_259 ( );
FILL FILL_24_DFFSR_259 ( );
FILL FILL_25_DFFSR_259 ( );
FILL FILL_26_DFFSR_259 ( );
FILL FILL_27_DFFSR_259 ( );
FILL FILL_28_DFFSR_259 ( );
FILL FILL_29_DFFSR_259 ( );
FILL FILL_30_DFFSR_259 ( );
FILL FILL_31_DFFSR_259 ( );
FILL FILL_32_DFFSR_259 ( );
FILL FILL_33_DFFSR_259 ( );
FILL FILL_34_DFFSR_259 ( );
FILL FILL_35_DFFSR_259 ( );
FILL FILL_36_DFFSR_259 ( );
FILL FILL_37_DFFSR_259 ( );
FILL FILL_38_DFFSR_259 ( );
FILL FILL_39_DFFSR_259 ( );
FILL FILL_40_DFFSR_259 ( );
FILL FILL_41_DFFSR_259 ( );
FILL FILL_42_DFFSR_259 ( );
FILL FILL_43_DFFSR_259 ( );
FILL FILL_44_DFFSR_259 ( );
FILL FILL_45_DFFSR_259 ( );
FILL FILL_46_DFFSR_259 ( );
FILL FILL_47_DFFSR_259 ( );
FILL FILL_48_DFFSR_259 ( );
FILL FILL_49_DFFSR_259 ( );
FILL FILL_50_DFFSR_259 ( );
FILL FILL_0_INVX1_183 ( );
FILL FILL_1_INVX1_183 ( );
FILL FILL_2_INVX1_183 ( );
FILL FILL_3_INVX1_183 ( );
FILL FILL_4_INVX1_183 ( );
FILL FILL_0_XOR2X1_7 ( );
FILL FILL_1_XOR2X1_7 ( );
FILL FILL_2_XOR2X1_7 ( );
FILL FILL_3_XOR2X1_7 ( );
FILL FILL_4_XOR2X1_7 ( );
FILL FILL_5_XOR2X1_7 ( );
FILL FILL_6_XOR2X1_7 ( );
FILL FILL_7_XOR2X1_7 ( );
FILL FILL_8_XOR2X1_7 ( );
FILL FILL_9_XOR2X1_7 ( );
FILL FILL_10_XOR2X1_7 ( );
FILL FILL_11_XOR2X1_7 ( );
FILL FILL_12_XOR2X1_7 ( );
FILL FILL_13_XOR2X1_7 ( );
FILL FILL_14_XOR2X1_7 ( );
FILL FILL_15_XOR2X1_7 ( );
FILL FILL_0_INVX1_171 ( );
FILL FILL_1_INVX1_171 ( );
FILL FILL_2_INVX1_171 ( );
FILL FILL_3_INVX1_171 ( );
FILL FILL_4_INVX1_171 ( );
FILL FILL_0_XNOR2X1_2 ( );
FILL FILL_1_XNOR2X1_2 ( );
FILL FILL_2_XNOR2X1_2 ( );
FILL FILL_3_XNOR2X1_2 ( );
FILL FILL_4_XNOR2X1_2 ( );
FILL FILL_5_XNOR2X1_2 ( );
FILL FILL_6_XNOR2X1_2 ( );
FILL FILL_7_XNOR2X1_2 ( );
FILL FILL_8_XNOR2X1_2 ( );
FILL FILL_9_XNOR2X1_2 ( );
FILL FILL_10_XNOR2X1_2 ( );
FILL FILL_11_XNOR2X1_2 ( );
FILL FILL_12_XNOR2X1_2 ( );
FILL FILL_13_XNOR2X1_2 ( );
FILL FILL_14_XNOR2X1_2 ( );
FILL FILL_15_XNOR2X1_2 ( );
FILL FILL_0_OAI21X1_84 ( );
FILL FILL_1_OAI21X1_84 ( );
FILL FILL_2_OAI21X1_84 ( );
FILL FILL_3_OAI21X1_84 ( );
FILL FILL_4_OAI21X1_84 ( );
FILL FILL_5_OAI21X1_84 ( );
FILL FILL_6_OAI21X1_84 ( );
FILL FILL_7_OAI21X1_84 ( );
FILL FILL_8_OAI21X1_84 ( );
FILL FILL_9_OAI21X1_84 ( );
FILL FILL_0_INVX1_180 ( );
FILL FILL_1_INVX1_180 ( );
FILL FILL_2_INVX1_180 ( );
FILL FILL_3_INVX1_180 ( );
FILL FILL_0_DFFSR_24 ( );
FILL FILL_1_DFFSR_24 ( );
FILL FILL_2_DFFSR_24 ( );
FILL FILL_3_DFFSR_24 ( );
FILL FILL_4_DFFSR_24 ( );
FILL FILL_5_DFFSR_24 ( );
FILL FILL_6_DFFSR_24 ( );
FILL FILL_7_DFFSR_24 ( );
FILL FILL_8_DFFSR_24 ( );
FILL FILL_9_DFFSR_24 ( );
FILL FILL_10_DFFSR_24 ( );
FILL FILL_11_DFFSR_24 ( );
FILL FILL_12_DFFSR_24 ( );
FILL FILL_13_DFFSR_24 ( );
FILL FILL_14_DFFSR_24 ( );
FILL FILL_15_DFFSR_24 ( );
FILL FILL_16_DFFSR_24 ( );
FILL FILL_17_DFFSR_24 ( );
FILL FILL_18_DFFSR_24 ( );
FILL FILL_19_DFFSR_24 ( );
FILL FILL_20_DFFSR_24 ( );
FILL FILL_21_DFFSR_24 ( );
FILL FILL_22_DFFSR_24 ( );
FILL FILL_23_DFFSR_24 ( );
FILL FILL_24_DFFSR_24 ( );
FILL FILL_25_DFFSR_24 ( );
FILL FILL_26_DFFSR_24 ( );
FILL FILL_27_DFFSR_24 ( );
FILL FILL_28_DFFSR_24 ( );
FILL FILL_29_DFFSR_24 ( );
FILL FILL_30_DFFSR_24 ( );
FILL FILL_31_DFFSR_24 ( );
FILL FILL_32_DFFSR_24 ( );
FILL FILL_33_DFFSR_24 ( );
FILL FILL_34_DFFSR_24 ( );
FILL FILL_35_DFFSR_24 ( );
FILL FILL_36_DFFSR_24 ( );
FILL FILL_37_DFFSR_24 ( );
FILL FILL_38_DFFSR_24 ( );
FILL FILL_39_DFFSR_24 ( );
FILL FILL_40_DFFSR_24 ( );
FILL FILL_41_DFFSR_24 ( );
FILL FILL_42_DFFSR_24 ( );
FILL FILL_43_DFFSR_24 ( );
FILL FILL_44_DFFSR_24 ( );
FILL FILL_45_DFFSR_24 ( );
FILL FILL_46_DFFSR_24 ( );
FILL FILL_47_DFFSR_24 ( );
FILL FILL_48_DFFSR_24 ( );
FILL FILL_49_DFFSR_24 ( );
FILL FILL_50_DFFSR_24 ( );
FILL FILL_51_DFFSR_24 ( );
FILL FILL_0_INVX1_56 ( );
FILL FILL_1_INVX1_56 ( );
FILL FILL_2_INVX1_56 ( );
FILL FILL_3_INVX1_56 ( );
FILL FILL_4_INVX1_56 ( );
FILL FILL_0_BUFX2_46 ( );
FILL FILL_1_BUFX2_46 ( );
FILL FILL_2_BUFX2_46 ( );
FILL FILL_3_BUFX2_46 ( );
FILL FILL_4_BUFX2_46 ( );
FILL FILL_5_BUFX2_46 ( );
FILL FILL_6_BUFX2_46 ( );
FILL FILL_0_DFFSR_38 ( );
FILL FILL_1_DFFSR_38 ( );
FILL FILL_2_DFFSR_38 ( );
FILL FILL_3_DFFSR_38 ( );
FILL FILL_4_DFFSR_38 ( );
FILL FILL_5_DFFSR_38 ( );
FILL FILL_6_DFFSR_38 ( );
FILL FILL_7_DFFSR_38 ( );
FILL FILL_8_DFFSR_38 ( );
FILL FILL_9_DFFSR_38 ( );
FILL FILL_10_DFFSR_38 ( );
FILL FILL_11_DFFSR_38 ( );
FILL FILL_12_DFFSR_38 ( );
FILL FILL_13_DFFSR_38 ( );
FILL FILL_14_DFFSR_38 ( );
FILL FILL_15_DFFSR_38 ( );
FILL FILL_16_DFFSR_38 ( );
FILL FILL_17_DFFSR_38 ( );
FILL FILL_18_DFFSR_38 ( );
FILL FILL_19_DFFSR_38 ( );
FILL FILL_20_DFFSR_38 ( );
FILL FILL_21_DFFSR_38 ( );
FILL FILL_22_DFFSR_38 ( );
FILL FILL_23_DFFSR_38 ( );
FILL FILL_24_DFFSR_38 ( );
FILL FILL_25_DFFSR_38 ( );
FILL FILL_26_DFFSR_38 ( );
FILL FILL_27_DFFSR_38 ( );
FILL FILL_28_DFFSR_38 ( );
FILL FILL_29_DFFSR_38 ( );
FILL FILL_30_DFFSR_38 ( );
FILL FILL_31_DFFSR_38 ( );
FILL FILL_32_DFFSR_38 ( );
FILL FILL_33_DFFSR_38 ( );
FILL FILL_34_DFFSR_38 ( );
FILL FILL_35_DFFSR_38 ( );
FILL FILL_36_DFFSR_38 ( );
FILL FILL_37_DFFSR_38 ( );
FILL FILL_38_DFFSR_38 ( );
FILL FILL_39_DFFSR_38 ( );
FILL FILL_40_DFFSR_38 ( );
FILL FILL_41_DFFSR_38 ( );
FILL FILL_42_DFFSR_38 ( );
FILL FILL_43_DFFSR_38 ( );
FILL FILL_44_DFFSR_38 ( );
FILL FILL_45_DFFSR_38 ( );
FILL FILL_46_DFFSR_38 ( );
FILL FILL_47_DFFSR_38 ( );
FILL FILL_48_DFFSR_38 ( );
FILL FILL_49_DFFSR_38 ( );
FILL FILL_50_DFFSR_38 ( );
FILL FILL_0_INVX1_14 ( );
FILL FILL_1_INVX1_14 ( );
FILL FILL_2_INVX1_14 ( );
FILL FILL_3_INVX1_14 ( );
FILL FILL_0_DFFSR_68 ( );
FILL FILL_1_DFFSR_68 ( );
FILL FILL_2_DFFSR_68 ( );
FILL FILL_3_DFFSR_68 ( );
FILL FILL_4_DFFSR_68 ( );
FILL FILL_5_DFFSR_68 ( );
FILL FILL_6_DFFSR_68 ( );
FILL FILL_7_DFFSR_68 ( );
FILL FILL_8_DFFSR_68 ( );
FILL FILL_9_DFFSR_68 ( );
FILL FILL_10_DFFSR_68 ( );
FILL FILL_11_DFFSR_68 ( );
FILL FILL_12_DFFSR_68 ( );
FILL FILL_13_DFFSR_68 ( );
FILL FILL_14_DFFSR_68 ( );
FILL FILL_15_DFFSR_68 ( );
FILL FILL_16_DFFSR_68 ( );
FILL FILL_17_DFFSR_68 ( );
FILL FILL_18_DFFSR_68 ( );
FILL FILL_19_DFFSR_68 ( );
FILL FILL_20_DFFSR_68 ( );
FILL FILL_21_DFFSR_68 ( );
FILL FILL_22_DFFSR_68 ( );
FILL FILL_23_DFFSR_68 ( );
FILL FILL_24_DFFSR_68 ( );
FILL FILL_25_DFFSR_68 ( );
FILL FILL_26_DFFSR_68 ( );
FILL FILL_27_DFFSR_68 ( );
FILL FILL_28_DFFSR_68 ( );
FILL FILL_29_DFFSR_68 ( );
FILL FILL_30_DFFSR_68 ( );
FILL FILL_31_DFFSR_68 ( );
FILL FILL_32_DFFSR_68 ( );
FILL FILL_33_DFFSR_68 ( );
FILL FILL_34_DFFSR_68 ( );
FILL FILL_35_DFFSR_68 ( );
FILL FILL_36_DFFSR_68 ( );
FILL FILL_37_DFFSR_68 ( );
FILL FILL_38_DFFSR_68 ( );
FILL FILL_39_DFFSR_68 ( );
FILL FILL_40_DFFSR_68 ( );
FILL FILL_41_DFFSR_68 ( );
FILL FILL_42_DFFSR_68 ( );
FILL FILL_43_DFFSR_68 ( );
FILL FILL_44_DFFSR_68 ( );
FILL FILL_45_DFFSR_68 ( );
FILL FILL_46_DFFSR_68 ( );
FILL FILL_47_DFFSR_68 ( );
FILL FILL_48_DFFSR_68 ( );
FILL FILL_49_DFFSR_68 ( );
FILL FILL_50_DFFSR_68 ( );
FILL FILL_0_NAND3X1_50 ( );
FILL FILL_1_NAND3X1_50 ( );
FILL FILL_2_NAND3X1_50 ( );
FILL FILL_3_NAND3X1_50 ( );
FILL FILL_4_NAND3X1_50 ( );
FILL FILL_5_NAND3X1_50 ( );
FILL FILL_6_NAND3X1_50 ( );
FILL FILL_7_NAND3X1_50 ( );
FILL FILL_8_NAND3X1_50 ( );
FILL FILL_0_INVX1_50 ( );
FILL FILL_1_INVX1_50 ( );
FILL FILL_2_INVX1_50 ( );
FILL FILL_3_INVX1_50 ( );
FILL FILL_4_INVX1_50 ( );
FILL FILL_0_NAND2X1_4 ( );
FILL FILL_1_NAND2X1_4 ( );
FILL FILL_2_NAND2X1_4 ( );
FILL FILL_3_NAND2X1_4 ( );
FILL FILL_4_NAND2X1_4 ( );
FILL FILL_5_NAND2X1_4 ( );
FILL FILL_6_NAND2X1_4 ( );
FILL FILL_0_NOR2X1_28 ( );
FILL FILL_1_NOR2X1_28 ( );
FILL FILL_2_NOR2X1_28 ( );
FILL FILL_3_NOR2X1_28 ( );
FILL FILL_4_NOR2X1_28 ( );
FILL FILL_5_NOR2X1_28 ( );
FILL FILL_6_NOR2X1_28 ( );
FILL FILL_0_INVX1_118 ( );
FILL FILL_1_INVX1_118 ( );
FILL FILL_2_INVX1_118 ( );
FILL FILL_3_INVX1_118 ( );
FILL FILL_4_INVX1_118 ( );
FILL FILL_0_XNOR2X1_4 ( );
FILL FILL_1_XNOR2X1_4 ( );
FILL FILL_2_XNOR2X1_4 ( );
FILL FILL_3_XNOR2X1_4 ( );
FILL FILL_4_XNOR2X1_4 ( );
FILL FILL_5_XNOR2X1_4 ( );
FILL FILL_6_XNOR2X1_4 ( );
FILL FILL_7_XNOR2X1_4 ( );
FILL FILL_8_XNOR2X1_4 ( );
FILL FILL_9_XNOR2X1_4 ( );
FILL FILL_10_XNOR2X1_4 ( );
FILL FILL_11_XNOR2X1_4 ( );
FILL FILL_12_XNOR2X1_4 ( );
FILL FILL_13_XNOR2X1_4 ( );
FILL FILL_14_XNOR2X1_4 ( );
FILL FILL_15_XNOR2X1_4 ( );
FILL FILL_0_DFFSR_43 ( );
FILL FILL_1_DFFSR_43 ( );
FILL FILL_2_DFFSR_43 ( );
FILL FILL_3_DFFSR_43 ( );
FILL FILL_4_DFFSR_43 ( );
FILL FILL_5_DFFSR_43 ( );
FILL FILL_6_DFFSR_43 ( );
FILL FILL_7_DFFSR_43 ( );
FILL FILL_8_DFFSR_43 ( );
FILL FILL_9_DFFSR_43 ( );
FILL FILL_10_DFFSR_43 ( );
FILL FILL_11_DFFSR_43 ( );
FILL FILL_12_DFFSR_43 ( );
FILL FILL_13_DFFSR_43 ( );
FILL FILL_14_DFFSR_43 ( );
FILL FILL_15_DFFSR_43 ( );
FILL FILL_16_DFFSR_43 ( );
FILL FILL_17_DFFSR_43 ( );
FILL FILL_18_DFFSR_43 ( );
FILL FILL_19_DFFSR_43 ( );
FILL FILL_20_DFFSR_43 ( );
FILL FILL_21_DFFSR_43 ( );
FILL FILL_22_DFFSR_43 ( );
FILL FILL_23_DFFSR_43 ( );
FILL FILL_24_DFFSR_43 ( );
FILL FILL_25_DFFSR_43 ( );
FILL FILL_26_DFFSR_43 ( );
FILL FILL_27_DFFSR_43 ( );
FILL FILL_28_DFFSR_43 ( );
FILL FILL_29_DFFSR_43 ( );
FILL FILL_30_DFFSR_43 ( );
FILL FILL_31_DFFSR_43 ( );
FILL FILL_32_DFFSR_43 ( );
FILL FILL_33_DFFSR_43 ( );
FILL FILL_34_DFFSR_43 ( );
FILL FILL_35_DFFSR_43 ( );
FILL FILL_36_DFFSR_43 ( );
FILL FILL_37_DFFSR_43 ( );
FILL FILL_38_DFFSR_43 ( );
FILL FILL_39_DFFSR_43 ( );
FILL FILL_40_DFFSR_43 ( );
FILL FILL_41_DFFSR_43 ( );
FILL FILL_42_DFFSR_43 ( );
FILL FILL_43_DFFSR_43 ( );
FILL FILL_44_DFFSR_43 ( );
FILL FILL_45_DFFSR_43 ( );
FILL FILL_46_DFFSR_43 ( );
FILL FILL_47_DFFSR_43 ( );
FILL FILL_48_DFFSR_43 ( );
FILL FILL_49_DFFSR_43 ( );
FILL FILL_50_DFFSR_43 ( );
FILL FILL_0_NAND3X1_1 ( );
FILL FILL_1_NAND3X1_1 ( );
FILL FILL_2_NAND3X1_1 ( );
FILL FILL_3_NAND3X1_1 ( );
FILL FILL_4_NAND3X1_1 ( );
FILL FILL_5_NAND3X1_1 ( );
FILL FILL_6_NAND3X1_1 ( );
FILL FILL_7_NAND3X1_1 ( );
FILL FILL_8_NAND3X1_1 ( );
FILL FILL_9_NAND3X1_1 ( );
FILL FILL_0_NOR2X1_6 ( );
FILL FILL_1_NOR2X1_6 ( );
FILL FILL_2_NOR2X1_6 ( );
FILL FILL_3_NOR2X1_6 ( );
FILL FILL_4_NOR2X1_6 ( );
FILL FILL_5_NOR2X1_6 ( );
FILL FILL_6_NOR2X1_6 ( );
FILL FILL_0_NAND2X1_11 ( );
FILL FILL_1_NAND2X1_11 ( );
FILL FILL_2_NAND2X1_11 ( );
FILL FILL_3_NAND2X1_11 ( );
FILL FILL_4_NAND2X1_11 ( );
FILL FILL_5_NAND2X1_11 ( );
FILL FILL_6_NAND2X1_11 ( );
FILL FILL_0_DFFSR_41 ( );
FILL FILL_1_DFFSR_41 ( );
FILL FILL_2_DFFSR_41 ( );
FILL FILL_3_DFFSR_41 ( );
FILL FILL_4_DFFSR_41 ( );
FILL FILL_5_DFFSR_41 ( );
FILL FILL_6_DFFSR_41 ( );
FILL FILL_7_DFFSR_41 ( );
FILL FILL_8_DFFSR_41 ( );
FILL FILL_9_DFFSR_41 ( );
FILL FILL_10_DFFSR_41 ( );
FILL FILL_11_DFFSR_41 ( );
FILL FILL_12_DFFSR_41 ( );
FILL FILL_13_DFFSR_41 ( );
FILL FILL_14_DFFSR_41 ( );
FILL FILL_15_DFFSR_41 ( );
FILL FILL_16_DFFSR_41 ( );
FILL FILL_17_DFFSR_41 ( );
FILL FILL_18_DFFSR_41 ( );
FILL FILL_19_DFFSR_41 ( );
FILL FILL_20_DFFSR_41 ( );
FILL FILL_21_DFFSR_41 ( );
FILL FILL_22_DFFSR_41 ( );
FILL FILL_23_DFFSR_41 ( );
FILL FILL_24_DFFSR_41 ( );
FILL FILL_25_DFFSR_41 ( );
FILL FILL_26_DFFSR_41 ( );
FILL FILL_27_DFFSR_41 ( );
FILL FILL_28_DFFSR_41 ( );
FILL FILL_29_DFFSR_41 ( );
FILL FILL_30_DFFSR_41 ( );
FILL FILL_31_DFFSR_41 ( );
FILL FILL_32_DFFSR_41 ( );
FILL FILL_33_DFFSR_41 ( );
FILL FILL_34_DFFSR_41 ( );
FILL FILL_35_DFFSR_41 ( );
FILL FILL_36_DFFSR_41 ( );
FILL FILL_37_DFFSR_41 ( );
FILL FILL_38_DFFSR_41 ( );
FILL FILL_39_DFFSR_41 ( );
FILL FILL_40_DFFSR_41 ( );
FILL FILL_41_DFFSR_41 ( );
FILL FILL_42_DFFSR_41 ( );
FILL FILL_43_DFFSR_41 ( );
FILL FILL_44_DFFSR_41 ( );
FILL FILL_45_DFFSR_41 ( );
FILL FILL_46_DFFSR_41 ( );
FILL FILL_47_DFFSR_41 ( );
FILL FILL_48_DFFSR_41 ( );
FILL FILL_49_DFFSR_41 ( );
FILL FILL_50_DFFSR_41 ( );
FILL FILL_0_CLKBUF1_3 ( );
FILL FILL_1_CLKBUF1_3 ( );
FILL FILL_2_CLKBUF1_3 ( );
FILL FILL_3_CLKBUF1_3 ( );
FILL FILL_4_CLKBUF1_3 ( );
FILL FILL_5_CLKBUF1_3 ( );
FILL FILL_6_CLKBUF1_3 ( );
FILL FILL_7_CLKBUF1_3 ( );
FILL FILL_8_CLKBUF1_3 ( );
FILL FILL_9_CLKBUF1_3 ( );
FILL FILL_10_CLKBUF1_3 ( );
FILL FILL_11_CLKBUF1_3 ( );
FILL FILL_12_CLKBUF1_3 ( );
FILL FILL_13_CLKBUF1_3 ( );
FILL FILL_14_CLKBUF1_3 ( );
FILL FILL_15_CLKBUF1_3 ( );
FILL FILL_16_CLKBUF1_3 ( );
FILL FILL_17_CLKBUF1_3 ( );
FILL FILL_18_CLKBUF1_3 ( );
FILL FILL_19_CLKBUF1_3 ( );
FILL FILL_20_CLKBUF1_3 ( );
FILL FILL_21_CLKBUF1_3 ( );
FILL FILL_0_NAND2X1_39 ( );
FILL FILL_1_NAND2X1_39 ( );
FILL FILL_2_NAND2X1_39 ( );
FILL FILL_3_NAND2X1_39 ( );
FILL FILL_4_NAND2X1_39 ( );
FILL FILL_5_NAND2X1_39 ( );
FILL FILL_6_NAND2X1_39 ( );
FILL FILL_0_INVX1_75 ( );
FILL FILL_1_INVX1_75 ( );
FILL FILL_2_INVX1_75 ( );
FILL FILL_3_INVX1_75 ( );
FILL FILL_4_INVX1_75 ( );
FILL FILL_0_DFFSR_210 ( );
FILL FILL_1_DFFSR_210 ( );
FILL FILL_2_DFFSR_210 ( );
FILL FILL_3_DFFSR_210 ( );
FILL FILL_4_DFFSR_210 ( );
FILL FILL_5_DFFSR_210 ( );
FILL FILL_6_DFFSR_210 ( );
FILL FILL_7_DFFSR_210 ( );
FILL FILL_8_DFFSR_210 ( );
FILL FILL_9_DFFSR_210 ( );
FILL FILL_10_DFFSR_210 ( );
FILL FILL_11_DFFSR_210 ( );
FILL FILL_12_DFFSR_210 ( );
FILL FILL_13_DFFSR_210 ( );
FILL FILL_14_DFFSR_210 ( );
FILL FILL_15_DFFSR_210 ( );
FILL FILL_16_DFFSR_210 ( );
FILL FILL_17_DFFSR_210 ( );
FILL FILL_18_DFFSR_210 ( );
FILL FILL_19_DFFSR_210 ( );
FILL FILL_20_DFFSR_210 ( );
FILL FILL_21_DFFSR_210 ( );
FILL FILL_22_DFFSR_210 ( );
FILL FILL_23_DFFSR_210 ( );
FILL FILL_24_DFFSR_210 ( );
FILL FILL_25_DFFSR_210 ( );
FILL FILL_26_DFFSR_210 ( );
FILL FILL_27_DFFSR_210 ( );
FILL FILL_28_DFFSR_210 ( );
FILL FILL_29_DFFSR_210 ( );
FILL FILL_30_DFFSR_210 ( );
FILL FILL_31_DFFSR_210 ( );
FILL FILL_32_DFFSR_210 ( );
FILL FILL_33_DFFSR_210 ( );
FILL FILL_34_DFFSR_210 ( );
FILL FILL_35_DFFSR_210 ( );
FILL FILL_36_DFFSR_210 ( );
FILL FILL_37_DFFSR_210 ( );
FILL FILL_38_DFFSR_210 ( );
FILL FILL_39_DFFSR_210 ( );
FILL FILL_40_DFFSR_210 ( );
FILL FILL_41_DFFSR_210 ( );
FILL FILL_42_DFFSR_210 ( );
FILL FILL_43_DFFSR_210 ( );
FILL FILL_44_DFFSR_210 ( );
FILL FILL_45_DFFSR_210 ( );
FILL FILL_46_DFFSR_210 ( );
FILL FILL_47_DFFSR_210 ( );
FILL FILL_48_DFFSR_210 ( );
FILL FILL_49_DFFSR_210 ( );
FILL FILL_50_DFFSR_210 ( );
FILL FILL_0_OAI21X1_90 ( );
FILL FILL_1_OAI21X1_90 ( );
FILL FILL_2_OAI21X1_90 ( );
FILL FILL_3_OAI21X1_90 ( );
FILL FILL_4_OAI21X1_90 ( );
FILL FILL_5_OAI21X1_90 ( );
FILL FILL_6_OAI21X1_90 ( );
FILL FILL_7_OAI21X1_90 ( );
FILL FILL_8_OAI21X1_90 ( );
FILL FILL_0_DFFSR_262 ( );
FILL FILL_1_DFFSR_262 ( );
FILL FILL_2_DFFSR_262 ( );
FILL FILL_3_DFFSR_262 ( );
FILL FILL_4_DFFSR_262 ( );
FILL FILL_5_DFFSR_262 ( );
FILL FILL_6_DFFSR_262 ( );
FILL FILL_7_DFFSR_262 ( );
FILL FILL_8_DFFSR_262 ( );
FILL FILL_9_DFFSR_262 ( );
FILL FILL_10_DFFSR_262 ( );
FILL FILL_11_DFFSR_262 ( );
FILL FILL_12_DFFSR_262 ( );
FILL FILL_13_DFFSR_262 ( );
FILL FILL_14_DFFSR_262 ( );
FILL FILL_15_DFFSR_262 ( );
FILL FILL_16_DFFSR_262 ( );
FILL FILL_17_DFFSR_262 ( );
FILL FILL_18_DFFSR_262 ( );
FILL FILL_19_DFFSR_262 ( );
FILL FILL_20_DFFSR_262 ( );
FILL FILL_21_DFFSR_262 ( );
FILL FILL_22_DFFSR_262 ( );
FILL FILL_23_DFFSR_262 ( );
FILL FILL_24_DFFSR_262 ( );
FILL FILL_25_DFFSR_262 ( );
FILL FILL_26_DFFSR_262 ( );
FILL FILL_27_DFFSR_262 ( );
FILL FILL_28_DFFSR_262 ( );
FILL FILL_29_DFFSR_262 ( );
FILL FILL_30_DFFSR_262 ( );
FILL FILL_31_DFFSR_262 ( );
FILL FILL_32_DFFSR_262 ( );
FILL FILL_33_DFFSR_262 ( );
FILL FILL_34_DFFSR_262 ( );
FILL FILL_35_DFFSR_262 ( );
FILL FILL_36_DFFSR_262 ( );
FILL FILL_37_DFFSR_262 ( );
FILL FILL_38_DFFSR_262 ( );
FILL FILL_39_DFFSR_262 ( );
FILL FILL_40_DFFSR_262 ( );
FILL FILL_41_DFFSR_262 ( );
FILL FILL_42_DFFSR_262 ( );
FILL FILL_43_DFFSR_262 ( );
FILL FILL_44_DFFSR_262 ( );
FILL FILL_45_DFFSR_262 ( );
FILL FILL_46_DFFSR_262 ( );
FILL FILL_47_DFFSR_262 ( );
FILL FILL_48_DFFSR_262 ( );
FILL FILL_49_DFFSR_262 ( );
FILL FILL_50_DFFSR_262 ( );
FILL FILL_0_CLKBUF1_47 ( );
FILL FILL_1_CLKBUF1_47 ( );
FILL FILL_2_CLKBUF1_47 ( );
FILL FILL_3_CLKBUF1_47 ( );
FILL FILL_4_CLKBUF1_47 ( );
FILL FILL_5_CLKBUF1_47 ( );
FILL FILL_6_CLKBUF1_47 ( );
FILL FILL_7_CLKBUF1_47 ( );
FILL FILL_8_CLKBUF1_47 ( );
FILL FILL_9_CLKBUF1_47 ( );
FILL FILL_10_CLKBUF1_47 ( );
FILL FILL_11_CLKBUF1_47 ( );
FILL FILL_12_CLKBUF1_47 ( );
FILL FILL_13_CLKBUF1_47 ( );
FILL FILL_14_CLKBUF1_47 ( );
FILL FILL_15_CLKBUF1_47 ( );
FILL FILL_16_CLKBUF1_47 ( );
FILL FILL_17_CLKBUF1_47 ( );
FILL FILL_18_CLKBUF1_47 ( );
FILL FILL_19_CLKBUF1_47 ( );
FILL FILL_20_CLKBUF1_47 ( );
FILL FILL_0_NAND2X1_153 ( );
FILL FILL_1_NAND2X1_153 ( );
FILL FILL_2_NAND2X1_153 ( );
FILL FILL_3_NAND2X1_153 ( );
FILL FILL_4_NAND2X1_153 ( );
FILL FILL_5_NAND2X1_153 ( );
FILL FILL_6_NAND2X1_153 ( );
FILL FILL_0_DFFSR_30 ( );
FILL FILL_1_DFFSR_30 ( );
FILL FILL_2_DFFSR_30 ( );
FILL FILL_3_DFFSR_30 ( );
FILL FILL_4_DFFSR_30 ( );
FILL FILL_5_DFFSR_30 ( );
FILL FILL_6_DFFSR_30 ( );
FILL FILL_7_DFFSR_30 ( );
FILL FILL_8_DFFSR_30 ( );
FILL FILL_9_DFFSR_30 ( );
FILL FILL_10_DFFSR_30 ( );
FILL FILL_11_DFFSR_30 ( );
FILL FILL_12_DFFSR_30 ( );
FILL FILL_13_DFFSR_30 ( );
FILL FILL_14_DFFSR_30 ( );
FILL FILL_15_DFFSR_30 ( );
FILL FILL_16_DFFSR_30 ( );
FILL FILL_17_DFFSR_30 ( );
FILL FILL_18_DFFSR_30 ( );
FILL FILL_19_DFFSR_30 ( );
FILL FILL_20_DFFSR_30 ( );
FILL FILL_21_DFFSR_30 ( );
FILL FILL_22_DFFSR_30 ( );
FILL FILL_23_DFFSR_30 ( );
FILL FILL_24_DFFSR_30 ( );
FILL FILL_25_DFFSR_30 ( );
FILL FILL_26_DFFSR_30 ( );
FILL FILL_27_DFFSR_30 ( );
FILL FILL_28_DFFSR_30 ( );
FILL FILL_29_DFFSR_30 ( );
FILL FILL_30_DFFSR_30 ( );
FILL FILL_31_DFFSR_30 ( );
FILL FILL_32_DFFSR_30 ( );
FILL FILL_33_DFFSR_30 ( );
FILL FILL_34_DFFSR_30 ( );
FILL FILL_35_DFFSR_30 ( );
FILL FILL_36_DFFSR_30 ( );
FILL FILL_37_DFFSR_30 ( );
FILL FILL_38_DFFSR_30 ( );
FILL FILL_39_DFFSR_30 ( );
FILL FILL_40_DFFSR_30 ( );
FILL FILL_41_DFFSR_30 ( );
FILL FILL_42_DFFSR_30 ( );
FILL FILL_43_DFFSR_30 ( );
FILL FILL_44_DFFSR_30 ( );
FILL FILL_45_DFFSR_30 ( );
FILL FILL_46_DFFSR_30 ( );
FILL FILL_47_DFFSR_30 ( );
FILL FILL_48_DFFSR_30 ( );
FILL FILL_49_DFFSR_30 ( );
FILL FILL_50_DFFSR_30 ( );
FILL FILL_51_DFFSR_30 ( );
FILL FILL_0_INVX1_57 ( );
FILL FILL_1_INVX1_57 ( );
FILL FILL_2_INVX1_57 ( );
FILL FILL_3_INVX1_57 ( );
FILL FILL_4_INVX1_57 ( );
FILL FILL_0_OAI22X1_24 ( );
FILL FILL_1_OAI22X1_24 ( );
FILL FILL_2_OAI22X1_24 ( );
FILL FILL_3_OAI22X1_24 ( );
FILL FILL_4_OAI22X1_24 ( );
FILL FILL_5_OAI22X1_24 ( );
FILL FILL_6_OAI22X1_24 ( );
FILL FILL_7_OAI22X1_24 ( );
FILL FILL_8_OAI22X1_24 ( );
FILL FILL_9_OAI22X1_24 ( );
FILL FILL_10_OAI22X1_24 ( );
FILL FILL_0_INVX1_15 ( );
FILL FILL_1_INVX1_15 ( );
FILL FILL_2_INVX1_15 ( );
FILL FILL_3_INVX1_15 ( );
FILL FILL_4_INVX1_15 ( );
FILL FILL_0_OAI22X1_6 ( );
FILL FILL_1_OAI22X1_6 ( );
FILL FILL_2_OAI22X1_6 ( );
FILL FILL_3_OAI22X1_6 ( );
FILL FILL_4_OAI22X1_6 ( );
FILL FILL_5_OAI22X1_6 ( );
FILL FILL_6_OAI22X1_6 ( );
FILL FILL_7_OAI22X1_6 ( );
FILL FILL_8_OAI22X1_6 ( );
FILL FILL_9_OAI22X1_6 ( );
FILL FILL_10_OAI22X1_6 ( );
FILL FILL_11_OAI22X1_6 ( );
FILL FILL_0_NAND2X1_14 ( );
FILL FILL_1_NAND2X1_14 ( );
FILL FILL_2_NAND2X1_14 ( );
FILL FILL_3_NAND2X1_14 ( );
FILL FILL_4_NAND2X1_14 ( );
FILL FILL_5_NAND2X1_14 ( );
FILL FILL_6_NAND2X1_14 ( );
FILL FILL_0_NOR2X1_7 ( );
FILL FILL_1_NOR2X1_7 ( );
FILL FILL_2_NOR2X1_7 ( );
FILL FILL_3_NOR2X1_7 ( );
FILL FILL_4_NOR2X1_7 ( );
FILL FILL_5_NOR2X1_7 ( );
FILL FILL_6_NOR2X1_7 ( );
FILL FILL_0_NAND2X1_6 ( );
FILL FILL_1_NAND2X1_6 ( );
FILL FILL_2_NAND2X1_6 ( );
FILL FILL_3_NAND2X1_6 ( );
FILL FILL_4_NAND2X1_6 ( );
FILL FILL_5_NAND2X1_6 ( );
FILL FILL_6_NAND2X1_6 ( );
FILL FILL_0_NOR2X1_10 ( );
FILL FILL_1_NOR2X1_10 ( );
FILL FILL_2_NOR2X1_10 ( );
FILL FILL_3_NOR2X1_10 ( );
FILL FILL_4_NOR2X1_10 ( );
FILL FILL_5_NOR2X1_10 ( );
FILL FILL_6_NOR2X1_10 ( );
FILL FILL_0_AND2X2_12 ( );
FILL FILL_1_AND2X2_12 ( );
FILL FILL_2_AND2X2_12 ( );
FILL FILL_3_AND2X2_12 ( );
FILL FILL_4_AND2X2_12 ( );
FILL FILL_5_AND2X2_12 ( );
FILL FILL_6_AND2X2_12 ( );
FILL FILL_7_AND2X2_12 ( );
FILL FILL_8_AND2X2_12 ( );
FILL FILL_0_OAI22X1_21 ( );
FILL FILL_1_OAI22X1_21 ( );
FILL FILL_2_OAI22X1_21 ( );
FILL FILL_3_OAI22X1_21 ( );
FILL FILL_4_OAI22X1_21 ( );
FILL FILL_5_OAI22X1_21 ( );
FILL FILL_6_OAI22X1_21 ( );
FILL FILL_7_OAI22X1_21 ( );
FILL FILL_8_OAI22X1_21 ( );
FILL FILL_9_OAI22X1_21 ( );
FILL FILL_10_OAI22X1_21 ( );
FILL FILL_11_OAI22X1_21 ( );
FILL FILL_0_BUFX2_18 ( );
FILL FILL_1_BUFX2_18 ( );
FILL FILL_2_BUFX2_18 ( );
FILL FILL_3_BUFX2_18 ( );
FILL FILL_4_BUFX2_18 ( );
FILL FILL_5_BUFX2_18 ( );
FILL FILL_6_BUFX2_18 ( );
FILL FILL_0_BUFX2_16 ( );
FILL FILL_1_BUFX2_16 ( );
FILL FILL_2_BUFX2_16 ( );
FILL FILL_3_BUFX2_16 ( );
FILL FILL_4_BUFX2_16 ( );
FILL FILL_5_BUFX2_16 ( );
FILL FILL_6_BUFX2_16 ( );
FILL FILL_0_AOI21X1_4 ( );
FILL FILL_1_AOI21X1_4 ( );
FILL FILL_2_AOI21X1_4 ( );
FILL FILL_3_AOI21X1_4 ( );
FILL FILL_4_AOI21X1_4 ( );
FILL FILL_5_AOI21X1_4 ( );
FILL FILL_6_AOI21X1_4 ( );
FILL FILL_7_AOI21X1_4 ( );
FILL FILL_8_AOI21X1_4 ( );
FILL FILL_9_AOI21X1_4 ( );
FILL FILL_0_OAI21X1_19 ( );
FILL FILL_1_OAI21X1_19 ( );
FILL FILL_2_OAI21X1_19 ( );
FILL FILL_3_OAI21X1_19 ( );
FILL FILL_4_OAI21X1_19 ( );
FILL FILL_5_OAI21X1_19 ( );
FILL FILL_6_OAI21X1_19 ( );
FILL FILL_7_OAI21X1_19 ( );
FILL FILL_8_OAI21X1_19 ( );
FILL FILL_0_DFFSR_69 ( );
FILL FILL_1_DFFSR_69 ( );
FILL FILL_2_DFFSR_69 ( );
FILL FILL_3_DFFSR_69 ( );
FILL FILL_4_DFFSR_69 ( );
FILL FILL_5_DFFSR_69 ( );
FILL FILL_6_DFFSR_69 ( );
FILL FILL_7_DFFSR_69 ( );
FILL FILL_8_DFFSR_69 ( );
FILL FILL_9_DFFSR_69 ( );
FILL FILL_10_DFFSR_69 ( );
FILL FILL_11_DFFSR_69 ( );
FILL FILL_12_DFFSR_69 ( );
FILL FILL_13_DFFSR_69 ( );
FILL FILL_14_DFFSR_69 ( );
FILL FILL_15_DFFSR_69 ( );
FILL FILL_16_DFFSR_69 ( );
FILL FILL_17_DFFSR_69 ( );
FILL FILL_18_DFFSR_69 ( );
FILL FILL_19_DFFSR_69 ( );
FILL FILL_20_DFFSR_69 ( );
FILL FILL_21_DFFSR_69 ( );
FILL FILL_22_DFFSR_69 ( );
FILL FILL_23_DFFSR_69 ( );
FILL FILL_24_DFFSR_69 ( );
FILL FILL_25_DFFSR_69 ( );
FILL FILL_26_DFFSR_69 ( );
FILL FILL_27_DFFSR_69 ( );
FILL FILL_28_DFFSR_69 ( );
FILL FILL_29_DFFSR_69 ( );
FILL FILL_30_DFFSR_69 ( );
FILL FILL_31_DFFSR_69 ( );
FILL FILL_32_DFFSR_69 ( );
FILL FILL_33_DFFSR_69 ( );
FILL FILL_34_DFFSR_69 ( );
FILL FILL_35_DFFSR_69 ( );
FILL FILL_36_DFFSR_69 ( );
FILL FILL_37_DFFSR_69 ( );
FILL FILL_38_DFFSR_69 ( );
FILL FILL_39_DFFSR_69 ( );
FILL FILL_40_DFFSR_69 ( );
FILL FILL_41_DFFSR_69 ( );
FILL FILL_42_DFFSR_69 ( );
FILL FILL_43_DFFSR_69 ( );
FILL FILL_44_DFFSR_69 ( );
FILL FILL_45_DFFSR_69 ( );
FILL FILL_46_DFFSR_69 ( );
FILL FILL_47_DFFSR_69 ( );
FILL FILL_48_DFFSR_69 ( );
FILL FILL_49_DFFSR_69 ( );
FILL FILL_50_DFFSR_69 ( );
FILL FILL_51_DFFSR_69 ( );
FILL FILL_0_NAND3X1_38 ( );
FILL FILL_1_NAND3X1_38 ( );
FILL FILL_2_NAND3X1_38 ( );
FILL FILL_3_NAND3X1_38 ( );
FILL FILL_4_NAND3X1_38 ( );
FILL FILL_5_NAND3X1_38 ( );
FILL FILL_6_NAND3X1_38 ( );
FILL FILL_7_NAND3X1_38 ( );
FILL FILL_8_NAND3X1_38 ( );
FILL FILL_9_NAND3X1_38 ( );
FILL FILL_0_DFFSR_77 ( );
FILL FILL_1_DFFSR_77 ( );
FILL FILL_2_DFFSR_77 ( );
FILL FILL_3_DFFSR_77 ( );
FILL FILL_4_DFFSR_77 ( );
FILL FILL_5_DFFSR_77 ( );
FILL FILL_6_DFFSR_77 ( );
FILL FILL_7_DFFSR_77 ( );
FILL FILL_8_DFFSR_77 ( );
FILL FILL_9_DFFSR_77 ( );
FILL FILL_10_DFFSR_77 ( );
FILL FILL_11_DFFSR_77 ( );
FILL FILL_12_DFFSR_77 ( );
FILL FILL_13_DFFSR_77 ( );
FILL FILL_14_DFFSR_77 ( );
FILL FILL_15_DFFSR_77 ( );
FILL FILL_16_DFFSR_77 ( );
FILL FILL_17_DFFSR_77 ( );
FILL FILL_18_DFFSR_77 ( );
FILL FILL_19_DFFSR_77 ( );
FILL FILL_20_DFFSR_77 ( );
FILL FILL_21_DFFSR_77 ( );
FILL FILL_22_DFFSR_77 ( );
FILL FILL_23_DFFSR_77 ( );
FILL FILL_24_DFFSR_77 ( );
FILL FILL_25_DFFSR_77 ( );
FILL FILL_26_DFFSR_77 ( );
FILL FILL_27_DFFSR_77 ( );
FILL FILL_28_DFFSR_77 ( );
FILL FILL_29_DFFSR_77 ( );
FILL FILL_30_DFFSR_77 ( );
FILL FILL_31_DFFSR_77 ( );
FILL FILL_32_DFFSR_77 ( );
FILL FILL_33_DFFSR_77 ( );
FILL FILL_34_DFFSR_77 ( );
FILL FILL_35_DFFSR_77 ( );
FILL FILL_36_DFFSR_77 ( );
FILL FILL_37_DFFSR_77 ( );
FILL FILL_38_DFFSR_77 ( );
FILL FILL_39_DFFSR_77 ( );
FILL FILL_40_DFFSR_77 ( );
FILL FILL_41_DFFSR_77 ( );
FILL FILL_42_DFFSR_77 ( );
FILL FILL_43_DFFSR_77 ( );
FILL FILL_44_DFFSR_77 ( );
FILL FILL_45_DFFSR_77 ( );
FILL FILL_46_DFFSR_77 ( );
FILL FILL_47_DFFSR_77 ( );
FILL FILL_48_DFFSR_77 ( );
FILL FILL_49_DFFSR_77 ( );
FILL FILL_50_DFFSR_77 ( );
FILL FILL_0_DFFSR_33 ( );
FILL FILL_1_DFFSR_33 ( );
FILL FILL_2_DFFSR_33 ( );
FILL FILL_3_DFFSR_33 ( );
FILL FILL_4_DFFSR_33 ( );
FILL FILL_5_DFFSR_33 ( );
FILL FILL_6_DFFSR_33 ( );
FILL FILL_7_DFFSR_33 ( );
FILL FILL_8_DFFSR_33 ( );
FILL FILL_9_DFFSR_33 ( );
FILL FILL_10_DFFSR_33 ( );
FILL FILL_11_DFFSR_33 ( );
FILL FILL_12_DFFSR_33 ( );
FILL FILL_13_DFFSR_33 ( );
FILL FILL_14_DFFSR_33 ( );
FILL FILL_15_DFFSR_33 ( );
FILL FILL_16_DFFSR_33 ( );
FILL FILL_17_DFFSR_33 ( );
FILL FILL_18_DFFSR_33 ( );
FILL FILL_19_DFFSR_33 ( );
FILL FILL_20_DFFSR_33 ( );
FILL FILL_21_DFFSR_33 ( );
FILL FILL_22_DFFSR_33 ( );
FILL FILL_23_DFFSR_33 ( );
FILL FILL_24_DFFSR_33 ( );
FILL FILL_25_DFFSR_33 ( );
FILL FILL_26_DFFSR_33 ( );
FILL FILL_27_DFFSR_33 ( );
FILL FILL_28_DFFSR_33 ( );
FILL FILL_29_DFFSR_33 ( );
FILL FILL_30_DFFSR_33 ( );
FILL FILL_31_DFFSR_33 ( );
FILL FILL_32_DFFSR_33 ( );
FILL FILL_33_DFFSR_33 ( );
FILL FILL_34_DFFSR_33 ( );
FILL FILL_35_DFFSR_33 ( );
FILL FILL_36_DFFSR_33 ( );
FILL FILL_37_DFFSR_33 ( );
FILL FILL_38_DFFSR_33 ( );
FILL FILL_39_DFFSR_33 ( );
FILL FILL_40_DFFSR_33 ( );
FILL FILL_41_DFFSR_33 ( );
FILL FILL_42_DFFSR_33 ( );
FILL FILL_43_DFFSR_33 ( );
FILL FILL_44_DFFSR_33 ( );
FILL FILL_45_DFFSR_33 ( );
FILL FILL_46_DFFSR_33 ( );
FILL FILL_47_DFFSR_33 ( );
FILL FILL_48_DFFSR_33 ( );
FILL FILL_49_DFFSR_33 ( );
FILL FILL_50_DFFSR_33 ( );
FILL FILL_51_DFFSR_33 ( );
FILL FILL_0_BUFX2_63 ( );
FILL FILL_1_BUFX2_63 ( );
FILL FILL_2_BUFX2_63 ( );
FILL FILL_3_BUFX2_63 ( );
FILL FILL_4_BUFX2_63 ( );
FILL FILL_5_BUFX2_63 ( );
FILL FILL_6_BUFX2_63 ( );
FILL FILL_0_DFFSR_218 ( );
FILL FILL_1_DFFSR_218 ( );
FILL FILL_2_DFFSR_218 ( );
FILL FILL_3_DFFSR_218 ( );
FILL FILL_4_DFFSR_218 ( );
FILL FILL_5_DFFSR_218 ( );
FILL FILL_6_DFFSR_218 ( );
FILL FILL_7_DFFSR_218 ( );
FILL FILL_8_DFFSR_218 ( );
FILL FILL_9_DFFSR_218 ( );
FILL FILL_10_DFFSR_218 ( );
FILL FILL_11_DFFSR_218 ( );
FILL FILL_12_DFFSR_218 ( );
FILL FILL_13_DFFSR_218 ( );
FILL FILL_14_DFFSR_218 ( );
FILL FILL_15_DFFSR_218 ( );
FILL FILL_16_DFFSR_218 ( );
FILL FILL_17_DFFSR_218 ( );
FILL FILL_18_DFFSR_218 ( );
FILL FILL_19_DFFSR_218 ( );
FILL FILL_20_DFFSR_218 ( );
FILL FILL_21_DFFSR_218 ( );
FILL FILL_22_DFFSR_218 ( );
FILL FILL_23_DFFSR_218 ( );
FILL FILL_24_DFFSR_218 ( );
FILL FILL_25_DFFSR_218 ( );
FILL FILL_26_DFFSR_218 ( );
FILL FILL_27_DFFSR_218 ( );
FILL FILL_28_DFFSR_218 ( );
FILL FILL_29_DFFSR_218 ( );
FILL FILL_30_DFFSR_218 ( );
FILL FILL_31_DFFSR_218 ( );
FILL FILL_32_DFFSR_218 ( );
FILL FILL_33_DFFSR_218 ( );
FILL FILL_34_DFFSR_218 ( );
FILL FILL_35_DFFSR_218 ( );
FILL FILL_36_DFFSR_218 ( );
FILL FILL_37_DFFSR_218 ( );
FILL FILL_38_DFFSR_218 ( );
FILL FILL_39_DFFSR_218 ( );
FILL FILL_40_DFFSR_218 ( );
FILL FILL_41_DFFSR_218 ( );
FILL FILL_42_DFFSR_218 ( );
FILL FILL_43_DFFSR_218 ( );
FILL FILL_44_DFFSR_218 ( );
FILL FILL_45_DFFSR_218 ( );
FILL FILL_46_DFFSR_218 ( );
FILL FILL_47_DFFSR_218 ( );
FILL FILL_48_DFFSR_218 ( );
FILL FILL_49_DFFSR_218 ( );
FILL FILL_50_DFFSR_218 ( );
FILL FILL_0_NAND2X1_121 ( );
FILL FILL_1_NAND2X1_121 ( );
FILL FILL_2_NAND2X1_121 ( );
FILL FILL_3_NAND2X1_121 ( );
FILL FILL_4_NAND2X1_121 ( );
FILL FILL_5_NAND2X1_121 ( );
FILL FILL_6_NAND2X1_121 ( );
FILL FILL_0_OR2X2_4 ( );
FILL FILL_1_OR2X2_4 ( );
FILL FILL_2_OR2X2_4 ( );
FILL FILL_3_OR2X2_4 ( );
FILL FILL_4_OR2X2_4 ( );
FILL FILL_5_OR2X2_4 ( );
FILL FILL_6_OR2X2_4 ( );
FILL FILL_7_OR2X2_4 ( );
FILL FILL_8_OR2X2_4 ( );
FILL FILL_0_AND2X2_40 ( );
FILL FILL_1_AND2X2_40 ( );
FILL FILL_2_AND2X2_40 ( );
FILL FILL_3_AND2X2_40 ( );
FILL FILL_4_AND2X2_40 ( );
FILL FILL_5_AND2X2_40 ( );
FILL FILL_6_AND2X2_40 ( );
FILL FILL_7_AND2X2_40 ( );
FILL FILL_8_AND2X2_40 ( );
FILL FILL_0_NAND2X1_114 ( );
FILL FILL_1_NAND2X1_114 ( );
FILL FILL_2_NAND2X1_114 ( );
FILL FILL_3_NAND2X1_114 ( );
FILL FILL_4_NAND2X1_114 ( );
FILL FILL_5_NAND2X1_114 ( );
FILL FILL_6_NAND2X1_114 ( );
FILL FILL_0_DFFSR_32 ( );
FILL FILL_1_DFFSR_32 ( );
FILL FILL_2_DFFSR_32 ( );
FILL FILL_3_DFFSR_32 ( );
FILL FILL_4_DFFSR_32 ( );
FILL FILL_5_DFFSR_32 ( );
FILL FILL_6_DFFSR_32 ( );
FILL FILL_7_DFFSR_32 ( );
FILL FILL_8_DFFSR_32 ( );
FILL FILL_9_DFFSR_32 ( );
FILL FILL_10_DFFSR_32 ( );
FILL FILL_11_DFFSR_32 ( );
FILL FILL_12_DFFSR_32 ( );
FILL FILL_13_DFFSR_32 ( );
FILL FILL_14_DFFSR_32 ( );
FILL FILL_15_DFFSR_32 ( );
FILL FILL_16_DFFSR_32 ( );
FILL FILL_17_DFFSR_32 ( );
FILL FILL_18_DFFSR_32 ( );
FILL FILL_19_DFFSR_32 ( );
FILL FILL_20_DFFSR_32 ( );
FILL FILL_21_DFFSR_32 ( );
FILL FILL_22_DFFSR_32 ( );
FILL FILL_23_DFFSR_32 ( );
FILL FILL_24_DFFSR_32 ( );
FILL FILL_25_DFFSR_32 ( );
FILL FILL_26_DFFSR_32 ( );
FILL FILL_27_DFFSR_32 ( );
FILL FILL_28_DFFSR_32 ( );
FILL FILL_29_DFFSR_32 ( );
FILL FILL_30_DFFSR_32 ( );
FILL FILL_31_DFFSR_32 ( );
FILL FILL_32_DFFSR_32 ( );
FILL FILL_33_DFFSR_32 ( );
FILL FILL_34_DFFSR_32 ( );
FILL FILL_35_DFFSR_32 ( );
FILL FILL_36_DFFSR_32 ( );
FILL FILL_37_DFFSR_32 ( );
FILL FILL_38_DFFSR_32 ( );
FILL FILL_39_DFFSR_32 ( );
FILL FILL_40_DFFSR_32 ( );
FILL FILL_41_DFFSR_32 ( );
FILL FILL_42_DFFSR_32 ( );
FILL FILL_43_DFFSR_32 ( );
FILL FILL_44_DFFSR_32 ( );
FILL FILL_45_DFFSR_32 ( );
FILL FILL_46_DFFSR_32 ( );
FILL FILL_47_DFFSR_32 ( );
FILL FILL_48_DFFSR_32 ( );
FILL FILL_49_DFFSR_32 ( );
FILL FILL_50_DFFSR_32 ( );
FILL FILL_0_DFFSR_22 ( );
FILL FILL_1_DFFSR_22 ( );
FILL FILL_2_DFFSR_22 ( );
FILL FILL_3_DFFSR_22 ( );
FILL FILL_4_DFFSR_22 ( );
FILL FILL_5_DFFSR_22 ( );
FILL FILL_6_DFFSR_22 ( );
FILL FILL_7_DFFSR_22 ( );
FILL FILL_8_DFFSR_22 ( );
FILL FILL_9_DFFSR_22 ( );
FILL FILL_10_DFFSR_22 ( );
FILL FILL_11_DFFSR_22 ( );
FILL FILL_12_DFFSR_22 ( );
FILL FILL_13_DFFSR_22 ( );
FILL FILL_14_DFFSR_22 ( );
FILL FILL_15_DFFSR_22 ( );
FILL FILL_16_DFFSR_22 ( );
FILL FILL_17_DFFSR_22 ( );
FILL FILL_18_DFFSR_22 ( );
FILL FILL_19_DFFSR_22 ( );
FILL FILL_20_DFFSR_22 ( );
FILL FILL_21_DFFSR_22 ( );
FILL FILL_22_DFFSR_22 ( );
FILL FILL_23_DFFSR_22 ( );
FILL FILL_24_DFFSR_22 ( );
FILL FILL_25_DFFSR_22 ( );
FILL FILL_26_DFFSR_22 ( );
FILL FILL_27_DFFSR_22 ( );
FILL FILL_28_DFFSR_22 ( );
FILL FILL_29_DFFSR_22 ( );
FILL FILL_30_DFFSR_22 ( );
FILL FILL_31_DFFSR_22 ( );
FILL FILL_32_DFFSR_22 ( );
FILL FILL_33_DFFSR_22 ( );
FILL FILL_34_DFFSR_22 ( );
FILL FILL_35_DFFSR_22 ( );
FILL FILL_36_DFFSR_22 ( );
FILL FILL_37_DFFSR_22 ( );
FILL FILL_38_DFFSR_22 ( );
FILL FILL_39_DFFSR_22 ( );
FILL FILL_40_DFFSR_22 ( );
FILL FILL_41_DFFSR_22 ( );
FILL FILL_42_DFFSR_22 ( );
FILL FILL_43_DFFSR_22 ( );
FILL FILL_44_DFFSR_22 ( );
FILL FILL_45_DFFSR_22 ( );
FILL FILL_46_DFFSR_22 ( );
FILL FILL_47_DFFSR_22 ( );
FILL FILL_48_DFFSR_22 ( );
FILL FILL_49_DFFSR_22 ( );
FILL FILL_50_DFFSR_22 ( );
FILL FILL_0_INVX1_42 ( );
FILL FILL_1_INVX1_42 ( );
FILL FILL_2_INVX1_42 ( );
FILL FILL_3_INVX1_42 ( );
FILL FILL_4_INVX1_42 ( );
FILL FILL_0_DFFSR_42 ( );
FILL FILL_1_DFFSR_42 ( );
FILL FILL_2_DFFSR_42 ( );
FILL FILL_3_DFFSR_42 ( );
FILL FILL_4_DFFSR_42 ( );
FILL FILL_5_DFFSR_42 ( );
FILL FILL_6_DFFSR_42 ( );
FILL FILL_7_DFFSR_42 ( );
FILL FILL_8_DFFSR_42 ( );
FILL FILL_9_DFFSR_42 ( );
FILL FILL_10_DFFSR_42 ( );
FILL FILL_11_DFFSR_42 ( );
FILL FILL_12_DFFSR_42 ( );
FILL FILL_13_DFFSR_42 ( );
FILL FILL_14_DFFSR_42 ( );
FILL FILL_15_DFFSR_42 ( );
FILL FILL_16_DFFSR_42 ( );
FILL FILL_17_DFFSR_42 ( );
FILL FILL_18_DFFSR_42 ( );
FILL FILL_19_DFFSR_42 ( );
FILL FILL_20_DFFSR_42 ( );
FILL FILL_21_DFFSR_42 ( );
FILL FILL_22_DFFSR_42 ( );
FILL FILL_23_DFFSR_42 ( );
FILL FILL_24_DFFSR_42 ( );
FILL FILL_25_DFFSR_42 ( );
FILL FILL_26_DFFSR_42 ( );
FILL FILL_27_DFFSR_42 ( );
FILL FILL_28_DFFSR_42 ( );
FILL FILL_29_DFFSR_42 ( );
FILL FILL_30_DFFSR_42 ( );
FILL FILL_31_DFFSR_42 ( );
FILL FILL_32_DFFSR_42 ( );
FILL FILL_33_DFFSR_42 ( );
FILL FILL_34_DFFSR_42 ( );
FILL FILL_35_DFFSR_42 ( );
FILL FILL_36_DFFSR_42 ( );
FILL FILL_37_DFFSR_42 ( );
FILL FILL_38_DFFSR_42 ( );
FILL FILL_39_DFFSR_42 ( );
FILL FILL_40_DFFSR_42 ( );
FILL FILL_41_DFFSR_42 ( );
FILL FILL_42_DFFSR_42 ( );
FILL FILL_43_DFFSR_42 ( );
FILL FILL_44_DFFSR_42 ( );
FILL FILL_45_DFFSR_42 ( );
FILL FILL_46_DFFSR_42 ( );
FILL FILL_47_DFFSR_42 ( );
FILL FILL_48_DFFSR_42 ( );
FILL FILL_49_DFFSR_42 ( );
FILL FILL_50_DFFSR_42 ( );
FILL FILL_51_DFFSR_42 ( );
FILL FILL_0_NAND3X1_29 ( );
FILL FILL_1_NAND3X1_29 ( );
FILL FILL_2_NAND3X1_29 ( );
FILL FILL_3_NAND3X1_29 ( );
FILL FILL_4_NAND3X1_29 ( );
FILL FILL_5_NAND3X1_29 ( );
FILL FILL_6_NAND3X1_29 ( );
FILL FILL_7_NAND3X1_29 ( );
FILL FILL_8_NAND3X1_29 ( );
FILL FILL_9_NAND3X1_29 ( );
FILL FILL_0_NAND3X1_12 ( );
FILL FILL_1_NAND3X1_12 ( );
FILL FILL_2_NAND3X1_12 ( );
FILL FILL_3_NAND3X1_12 ( );
FILL FILL_4_NAND3X1_12 ( );
FILL FILL_5_NAND3X1_12 ( );
FILL FILL_6_NAND3X1_12 ( );
FILL FILL_7_NAND3X1_12 ( );
FILL FILL_8_NAND3X1_12 ( );
FILL FILL_0_AND2X2_7 ( );
FILL FILL_1_AND2X2_7 ( );
FILL FILL_2_AND2X2_7 ( );
FILL FILL_3_AND2X2_7 ( );
FILL FILL_4_AND2X2_7 ( );
FILL FILL_5_AND2X2_7 ( );
FILL FILL_6_AND2X2_7 ( );
FILL FILL_7_AND2X2_7 ( );
FILL FILL_8_AND2X2_7 ( );
FILL FILL_0_NAND3X1_59 ( );
FILL FILL_1_NAND3X1_59 ( );
FILL FILL_2_NAND3X1_59 ( );
FILL FILL_3_NAND3X1_59 ( );
FILL FILL_4_NAND3X1_59 ( );
FILL FILL_5_NAND3X1_59 ( );
FILL FILL_6_NAND3X1_59 ( );
FILL FILL_7_NAND3X1_59 ( );
FILL FILL_8_NAND3X1_59 ( );
FILL FILL_0_BUFX2_1 ( );
FILL FILL_1_BUFX2_1 ( );
FILL FILL_2_BUFX2_1 ( );
FILL FILL_3_BUFX2_1 ( );
FILL FILL_4_BUFX2_1 ( );
FILL FILL_5_BUFX2_1 ( );
FILL FILL_6_BUFX2_1 ( );
FILL FILL_0_BUFX2_21 ( );
FILL FILL_1_BUFX2_21 ( );
FILL FILL_2_BUFX2_21 ( );
FILL FILL_3_BUFX2_21 ( );
FILL FILL_4_BUFX2_21 ( );
FILL FILL_5_BUFX2_21 ( );
FILL FILL_6_BUFX2_21 ( );
FILL FILL_0_NAND3X1_11 ( );
FILL FILL_1_NAND3X1_11 ( );
FILL FILL_2_NAND3X1_11 ( );
FILL FILL_3_NAND3X1_11 ( );
FILL FILL_4_NAND3X1_11 ( );
FILL FILL_5_NAND3X1_11 ( );
FILL FILL_6_NAND3X1_11 ( );
FILL FILL_7_NAND3X1_11 ( );
FILL FILL_8_NAND3X1_11 ( );
FILL FILL_9_NAND3X1_11 ( );
FILL FILL_0_NAND3X1_64 ( );
FILL FILL_1_NAND3X1_64 ( );
FILL FILL_2_NAND3X1_64 ( );
FILL FILL_3_NAND3X1_64 ( );
FILL FILL_4_NAND3X1_64 ( );
FILL FILL_5_NAND3X1_64 ( );
FILL FILL_6_NAND3X1_64 ( );
FILL FILL_7_NAND3X1_64 ( );
FILL FILL_8_NAND3X1_64 ( );
FILL FILL_0_BUFX2_14 ( );
FILL FILL_1_BUFX2_14 ( );
FILL FILL_2_BUFX2_14 ( );
FILL FILL_3_BUFX2_14 ( );
FILL FILL_4_BUFX2_14 ( );
FILL FILL_5_BUFX2_14 ( );
FILL FILL_6_BUFX2_14 ( );
FILL FILL_0_DFFPOSX1_8 ( );
FILL FILL_1_DFFPOSX1_8 ( );
FILL FILL_2_DFFPOSX1_8 ( );
FILL FILL_3_DFFPOSX1_8 ( );
FILL FILL_4_DFFPOSX1_8 ( );
FILL FILL_5_DFFPOSX1_8 ( );
FILL FILL_6_DFFPOSX1_8 ( );
FILL FILL_7_DFFPOSX1_8 ( );
FILL FILL_8_DFFPOSX1_8 ( );
FILL FILL_9_DFFPOSX1_8 ( );
FILL FILL_10_DFFPOSX1_8 ( );
FILL FILL_11_DFFPOSX1_8 ( );
FILL FILL_12_DFFPOSX1_8 ( );
FILL FILL_13_DFFPOSX1_8 ( );
FILL FILL_14_DFFPOSX1_8 ( );
FILL FILL_15_DFFPOSX1_8 ( );
FILL FILL_16_DFFPOSX1_8 ( );
FILL FILL_17_DFFPOSX1_8 ( );
FILL FILL_18_DFFPOSX1_8 ( );
FILL FILL_19_DFFPOSX1_8 ( );
FILL FILL_20_DFFPOSX1_8 ( );
FILL FILL_21_DFFPOSX1_8 ( );
FILL FILL_22_DFFPOSX1_8 ( );
FILL FILL_23_DFFPOSX1_8 ( );
FILL FILL_24_DFFPOSX1_8 ( );
FILL FILL_25_DFFPOSX1_8 ( );
FILL FILL_26_DFFPOSX1_8 ( );
FILL FILL_27_DFFPOSX1_8 ( );
FILL FILL_0_BUFX2_20 ( );
FILL FILL_1_BUFX2_20 ( );
FILL FILL_2_BUFX2_20 ( );
FILL FILL_3_BUFX2_20 ( );
FILL FILL_4_BUFX2_20 ( );
FILL FILL_5_BUFX2_20 ( );
FILL FILL_6_BUFX2_20 ( );
FILL FILL_0_NAND3X1_37 ( );
FILL FILL_1_NAND3X1_37 ( );
FILL FILL_2_NAND3X1_37 ( );
FILL FILL_3_NAND3X1_37 ( );
FILL FILL_4_NAND3X1_37 ( );
FILL FILL_5_NAND3X1_37 ( );
FILL FILL_6_NAND3X1_37 ( );
FILL FILL_7_NAND3X1_37 ( );
FILL FILL_8_NAND3X1_37 ( );
FILL FILL_0_NAND3X1_39 ( );
FILL FILL_1_NAND3X1_39 ( );
FILL FILL_2_NAND3X1_39 ( );
FILL FILL_3_NAND3X1_39 ( );
FILL FILL_4_NAND3X1_39 ( );
FILL FILL_5_NAND3X1_39 ( );
FILL FILL_6_NAND3X1_39 ( );
FILL FILL_7_NAND3X1_39 ( );
FILL FILL_8_NAND3X1_39 ( );
FILL FILL_9_NAND3X1_39 ( );
FILL FILL_0_NOR2X1_20 ( );
FILL FILL_1_NOR2X1_20 ( );
FILL FILL_2_NOR2X1_20 ( );
FILL FILL_3_NOR2X1_20 ( );
FILL FILL_4_NOR2X1_20 ( );
FILL FILL_5_NOR2X1_20 ( );
FILL FILL_6_NOR2X1_20 ( );
FILL FILL_0_INVX1_21 ( );
FILL FILL_1_INVX1_21 ( );
FILL FILL_2_INVX1_21 ( );
FILL FILL_3_INVX1_21 ( );
FILL FILL_4_INVX1_21 ( );
FILL FILL_0_DFFSR_112 ( );
FILL FILL_1_DFFSR_112 ( );
FILL FILL_2_DFFSR_112 ( );
FILL FILL_3_DFFSR_112 ( );
FILL FILL_4_DFFSR_112 ( );
FILL FILL_5_DFFSR_112 ( );
FILL FILL_6_DFFSR_112 ( );
FILL FILL_7_DFFSR_112 ( );
FILL FILL_8_DFFSR_112 ( );
FILL FILL_9_DFFSR_112 ( );
FILL FILL_10_DFFSR_112 ( );
FILL FILL_11_DFFSR_112 ( );
FILL FILL_12_DFFSR_112 ( );
FILL FILL_13_DFFSR_112 ( );
FILL FILL_14_DFFSR_112 ( );
FILL FILL_15_DFFSR_112 ( );
FILL FILL_16_DFFSR_112 ( );
FILL FILL_17_DFFSR_112 ( );
FILL FILL_18_DFFSR_112 ( );
FILL FILL_19_DFFSR_112 ( );
FILL FILL_20_DFFSR_112 ( );
FILL FILL_21_DFFSR_112 ( );
FILL FILL_22_DFFSR_112 ( );
FILL FILL_23_DFFSR_112 ( );
FILL FILL_24_DFFSR_112 ( );
FILL FILL_25_DFFSR_112 ( );
FILL FILL_26_DFFSR_112 ( );
FILL FILL_27_DFFSR_112 ( );
FILL FILL_28_DFFSR_112 ( );
FILL FILL_29_DFFSR_112 ( );
FILL FILL_30_DFFSR_112 ( );
FILL FILL_31_DFFSR_112 ( );
FILL FILL_32_DFFSR_112 ( );
FILL FILL_33_DFFSR_112 ( );
FILL FILL_34_DFFSR_112 ( );
FILL FILL_35_DFFSR_112 ( );
FILL FILL_36_DFFSR_112 ( );
FILL FILL_37_DFFSR_112 ( );
FILL FILL_38_DFFSR_112 ( );
FILL FILL_39_DFFSR_112 ( );
FILL FILL_40_DFFSR_112 ( );
FILL FILL_41_DFFSR_112 ( );
FILL FILL_42_DFFSR_112 ( );
FILL FILL_43_DFFSR_112 ( );
FILL FILL_44_DFFSR_112 ( );
FILL FILL_45_DFFSR_112 ( );
FILL FILL_46_DFFSR_112 ( );
FILL FILL_47_DFFSR_112 ( );
FILL FILL_48_DFFSR_112 ( );
FILL FILL_49_DFFSR_112 ( );
FILL FILL_50_DFFSR_112 ( );
FILL FILL_0_BUFX2_2 ( );
FILL FILL_1_BUFX2_2 ( );
FILL FILL_2_BUFX2_2 ( );
FILL FILL_3_BUFX2_2 ( );
FILL FILL_4_BUFX2_2 ( );
FILL FILL_5_BUFX2_2 ( );
FILL FILL_6_BUFX2_2 ( );
FILL FILL_0_INVX1_7 ( );
FILL FILL_1_INVX1_7 ( );
FILL FILL_2_INVX1_7 ( );
FILL FILL_3_INVX1_7 ( );
FILL FILL_4_INVX1_7 ( );
FILL FILL_0_INVX1_22 ( );
FILL FILL_1_INVX1_22 ( );
FILL FILL_2_INVX1_22 ( );
FILL FILL_3_INVX1_22 ( );
FILL FILL_0_CLKBUF1_7 ( );
FILL FILL_1_CLKBUF1_7 ( );
FILL FILL_2_CLKBUF1_7 ( );
FILL FILL_3_CLKBUF1_7 ( );
FILL FILL_4_CLKBUF1_7 ( );
FILL FILL_5_CLKBUF1_7 ( );
FILL FILL_6_CLKBUF1_7 ( );
FILL FILL_7_CLKBUF1_7 ( );
FILL FILL_8_CLKBUF1_7 ( );
FILL FILL_9_CLKBUF1_7 ( );
FILL FILL_10_CLKBUF1_7 ( );
FILL FILL_11_CLKBUF1_7 ( );
FILL FILL_12_CLKBUF1_7 ( );
FILL FILL_13_CLKBUF1_7 ( );
FILL FILL_14_CLKBUF1_7 ( );
FILL FILL_15_CLKBUF1_7 ( );
FILL FILL_16_CLKBUF1_7 ( );
FILL FILL_17_CLKBUF1_7 ( );
FILL FILL_18_CLKBUF1_7 ( );
FILL FILL_19_CLKBUF1_7 ( );
FILL FILL_20_CLKBUF1_7 ( );
FILL FILL_0_BUFX2_96 ( );
FILL FILL_1_BUFX2_96 ( );
FILL FILL_2_BUFX2_96 ( );
FILL FILL_3_BUFX2_96 ( );
FILL FILL_4_BUFX2_96 ( );
FILL FILL_5_BUFX2_96 ( );
FILL FILL_6_BUFX2_96 ( );
FILL FILL_0_DFFSR_255 ( );
FILL FILL_1_DFFSR_255 ( );
FILL FILL_2_DFFSR_255 ( );
FILL FILL_3_DFFSR_255 ( );
FILL FILL_4_DFFSR_255 ( );
FILL FILL_5_DFFSR_255 ( );
FILL FILL_6_DFFSR_255 ( );
FILL FILL_7_DFFSR_255 ( );
FILL FILL_8_DFFSR_255 ( );
FILL FILL_9_DFFSR_255 ( );
FILL FILL_10_DFFSR_255 ( );
FILL FILL_11_DFFSR_255 ( );
FILL FILL_12_DFFSR_255 ( );
FILL FILL_13_DFFSR_255 ( );
FILL FILL_14_DFFSR_255 ( );
FILL FILL_15_DFFSR_255 ( );
FILL FILL_16_DFFSR_255 ( );
FILL FILL_17_DFFSR_255 ( );
FILL FILL_18_DFFSR_255 ( );
FILL FILL_19_DFFSR_255 ( );
FILL FILL_20_DFFSR_255 ( );
FILL FILL_21_DFFSR_255 ( );
FILL FILL_22_DFFSR_255 ( );
FILL FILL_23_DFFSR_255 ( );
FILL FILL_24_DFFSR_255 ( );
FILL FILL_25_DFFSR_255 ( );
FILL FILL_26_DFFSR_255 ( );
FILL FILL_27_DFFSR_255 ( );
FILL FILL_28_DFFSR_255 ( );
FILL FILL_29_DFFSR_255 ( );
FILL FILL_30_DFFSR_255 ( );
FILL FILL_31_DFFSR_255 ( );
FILL FILL_32_DFFSR_255 ( );
FILL FILL_33_DFFSR_255 ( );
FILL FILL_34_DFFSR_255 ( );
FILL FILL_35_DFFSR_255 ( );
FILL FILL_36_DFFSR_255 ( );
FILL FILL_37_DFFSR_255 ( );
FILL FILL_38_DFFSR_255 ( );
FILL FILL_39_DFFSR_255 ( );
FILL FILL_40_DFFSR_255 ( );
FILL FILL_41_DFFSR_255 ( );
FILL FILL_42_DFFSR_255 ( );
FILL FILL_43_DFFSR_255 ( );
FILL FILL_44_DFFSR_255 ( );
FILL FILL_45_DFFSR_255 ( );
FILL FILL_46_DFFSR_255 ( );
FILL FILL_47_DFFSR_255 ( );
FILL FILL_48_DFFSR_255 ( );
FILL FILL_49_DFFSR_255 ( );
FILL FILL_50_DFFSR_255 ( );
FILL FILL_0_XOR2X1_8 ( );
FILL FILL_1_XOR2X1_8 ( );
FILL FILL_2_XOR2X1_8 ( );
FILL FILL_3_XOR2X1_8 ( );
FILL FILL_4_XOR2X1_8 ( );
FILL FILL_5_XOR2X1_8 ( );
FILL FILL_6_XOR2X1_8 ( );
FILL FILL_7_XOR2X1_8 ( );
FILL FILL_8_XOR2X1_8 ( );
FILL FILL_9_XOR2X1_8 ( );
FILL FILL_10_XOR2X1_8 ( );
FILL FILL_11_XOR2X1_8 ( );
FILL FILL_12_XOR2X1_8 ( );
FILL FILL_13_XOR2X1_8 ( );
FILL FILL_14_XOR2X1_8 ( );
FILL FILL_15_XOR2X1_8 ( );
FILL FILL_0_NAND2X1_112 ( );
FILL FILL_1_NAND2X1_112 ( );
FILL FILL_2_NAND2X1_112 ( );
FILL FILL_3_NAND2X1_112 ( );
FILL FILL_4_NAND2X1_112 ( );
FILL FILL_5_NAND2X1_112 ( );
FILL FILL_6_NAND2X1_112 ( );
FILL FILL_0_INVX1_174 ( );
FILL FILL_1_INVX1_174 ( );
FILL FILL_2_INVX1_174 ( );
FILL FILL_3_INVX1_174 ( );
FILL FILL_4_INVX1_174 ( );
FILL FILL_0_NAND3X1_245 ( );
FILL FILL_1_NAND3X1_245 ( );
FILL FILL_2_NAND3X1_245 ( );
FILL FILL_3_NAND3X1_245 ( );
FILL FILL_4_NAND3X1_245 ( );
FILL FILL_5_NAND3X1_245 ( );
FILL FILL_6_NAND3X1_245 ( );
FILL FILL_7_NAND3X1_245 ( );
FILL FILL_8_NAND3X1_245 ( );
FILL FILL_9_NAND3X1_245 ( );
FILL FILL_0_NAND2X1_113 ( );
FILL FILL_1_NAND2X1_113 ( );
FILL FILL_2_NAND2X1_113 ( );
FILL FILL_3_NAND2X1_113 ( );
FILL FILL_4_NAND2X1_113 ( );
FILL FILL_5_NAND2X1_113 ( );
FILL FILL_6_NAND2X1_113 ( );
FILL FILL_0_NAND3X1_246 ( );
FILL FILL_1_NAND3X1_246 ( );
FILL FILL_2_NAND3X1_246 ( );
FILL FILL_3_NAND3X1_246 ( );
FILL FILL_4_NAND3X1_246 ( );
FILL FILL_5_NAND3X1_246 ( );
FILL FILL_6_NAND3X1_246 ( );
FILL FILL_7_NAND3X1_246 ( );
FILL FILL_8_NAND3X1_246 ( );
FILL FILL_0_CLKBUF1_28 ( );
FILL FILL_1_CLKBUF1_28 ( );
FILL FILL_2_CLKBUF1_28 ( );
FILL FILL_3_CLKBUF1_28 ( );
FILL FILL_4_CLKBUF1_28 ( );
FILL FILL_5_CLKBUF1_28 ( );
FILL FILL_6_CLKBUF1_28 ( );
FILL FILL_7_CLKBUF1_28 ( );
FILL FILL_8_CLKBUF1_28 ( );
FILL FILL_9_CLKBUF1_28 ( );
FILL FILL_10_CLKBUF1_28 ( );
FILL FILL_11_CLKBUF1_28 ( );
FILL FILL_12_CLKBUF1_28 ( );
FILL FILL_13_CLKBUF1_28 ( );
FILL FILL_14_CLKBUF1_28 ( );
FILL FILL_15_CLKBUF1_28 ( );
FILL FILL_16_CLKBUF1_28 ( );
FILL FILL_17_CLKBUF1_28 ( );
FILL FILL_18_CLKBUF1_28 ( );
FILL FILL_19_CLKBUF1_28 ( );
FILL FILL_20_CLKBUF1_28 ( );
FILL FILL_0_NAND2X1_154 ( );
FILL FILL_1_NAND2X1_154 ( );
FILL FILL_2_NAND2X1_154 ( );
FILL FILL_3_NAND2X1_154 ( );
FILL FILL_4_NAND2X1_154 ( );
FILL FILL_5_NAND2X1_154 ( );
FILL FILL_6_NAND2X1_154 ( );
FILL FILL_0_DFFSR_40 ( );
FILL FILL_1_DFFSR_40 ( );
FILL FILL_2_DFFSR_40 ( );
FILL FILL_3_DFFSR_40 ( );
FILL FILL_4_DFFSR_40 ( );
FILL FILL_5_DFFSR_40 ( );
FILL FILL_6_DFFSR_40 ( );
FILL FILL_7_DFFSR_40 ( );
FILL FILL_8_DFFSR_40 ( );
FILL FILL_9_DFFSR_40 ( );
FILL FILL_10_DFFSR_40 ( );
FILL FILL_11_DFFSR_40 ( );
FILL FILL_12_DFFSR_40 ( );
FILL FILL_13_DFFSR_40 ( );
FILL FILL_14_DFFSR_40 ( );
FILL FILL_15_DFFSR_40 ( );
FILL FILL_16_DFFSR_40 ( );
FILL FILL_17_DFFSR_40 ( );
FILL FILL_18_DFFSR_40 ( );
FILL FILL_19_DFFSR_40 ( );
FILL FILL_20_DFFSR_40 ( );
FILL FILL_21_DFFSR_40 ( );
FILL FILL_22_DFFSR_40 ( );
FILL FILL_23_DFFSR_40 ( );
FILL FILL_24_DFFSR_40 ( );
FILL FILL_25_DFFSR_40 ( );
FILL FILL_26_DFFSR_40 ( );
FILL FILL_27_DFFSR_40 ( );
FILL FILL_28_DFFSR_40 ( );
FILL FILL_29_DFFSR_40 ( );
FILL FILL_30_DFFSR_40 ( );
FILL FILL_31_DFFSR_40 ( );
FILL FILL_32_DFFSR_40 ( );
FILL FILL_33_DFFSR_40 ( );
FILL FILL_34_DFFSR_40 ( );
FILL FILL_35_DFFSR_40 ( );
FILL FILL_36_DFFSR_40 ( );
FILL FILL_37_DFFSR_40 ( );
FILL FILL_38_DFFSR_40 ( );
FILL FILL_39_DFFSR_40 ( );
FILL FILL_40_DFFSR_40 ( );
FILL FILL_41_DFFSR_40 ( );
FILL FILL_42_DFFSR_40 ( );
FILL FILL_43_DFFSR_40 ( );
FILL FILL_44_DFFSR_40 ( );
FILL FILL_45_DFFSR_40 ( );
FILL FILL_46_DFFSR_40 ( );
FILL FILL_47_DFFSR_40 ( );
FILL FILL_48_DFFSR_40 ( );
FILL FILL_49_DFFSR_40 ( );
FILL FILL_50_DFFSR_40 ( );
FILL FILL_0_INVX1_43 ( );
FILL FILL_1_INVX1_43 ( );
FILL FILL_2_INVX1_43 ( );
FILL FILL_3_INVX1_43 ( );
FILL FILL_0_OAI22X1_18 ( );
FILL FILL_1_OAI22X1_18 ( );
FILL FILL_2_OAI22X1_18 ( );
FILL FILL_3_OAI22X1_18 ( );
FILL FILL_4_OAI22X1_18 ( );
FILL FILL_5_OAI22X1_18 ( );
FILL FILL_6_OAI22X1_18 ( );
FILL FILL_7_OAI22X1_18 ( );
FILL FILL_8_OAI22X1_18 ( );
FILL FILL_9_OAI22X1_18 ( );
FILL FILL_10_OAI22X1_18 ( );
FILL FILL_11_OAI22X1_18 ( );
FILL FILL_0_CLKBUF1_41 ( );
FILL FILL_1_CLKBUF1_41 ( );
FILL FILL_2_CLKBUF1_41 ( );
FILL FILL_3_CLKBUF1_41 ( );
FILL FILL_4_CLKBUF1_41 ( );
FILL FILL_5_CLKBUF1_41 ( );
FILL FILL_6_CLKBUF1_41 ( );
FILL FILL_7_CLKBUF1_41 ( );
FILL FILL_8_CLKBUF1_41 ( );
FILL FILL_9_CLKBUF1_41 ( );
FILL FILL_10_CLKBUF1_41 ( );
FILL FILL_11_CLKBUF1_41 ( );
FILL FILL_12_CLKBUF1_41 ( );
FILL FILL_13_CLKBUF1_41 ( );
FILL FILL_14_CLKBUF1_41 ( );
FILL FILL_15_CLKBUF1_41 ( );
FILL FILL_16_CLKBUF1_41 ( );
FILL FILL_17_CLKBUF1_41 ( );
FILL FILL_18_CLKBUF1_41 ( );
FILL FILL_19_CLKBUF1_41 ( );
FILL FILL_20_CLKBUF1_41 ( );
FILL FILL_0_NAND2X1_5 ( );
FILL FILL_1_NAND2X1_5 ( );
FILL FILL_2_NAND2X1_5 ( );
FILL FILL_3_NAND2X1_5 ( );
FILL FILL_4_NAND2X1_5 ( );
FILL FILL_5_NAND2X1_5 ( );
FILL FILL_6_NAND2X1_5 ( );
FILL FILL_0_NAND3X1_9 ( );
FILL FILL_1_NAND3X1_9 ( );
FILL FILL_2_NAND3X1_9 ( );
FILL FILL_3_NAND3X1_9 ( );
FILL FILL_4_NAND3X1_9 ( );
FILL FILL_5_NAND3X1_9 ( );
FILL FILL_6_NAND3X1_9 ( );
FILL FILL_7_NAND3X1_9 ( );
FILL FILL_8_NAND3X1_9 ( );
FILL FILL_0_NAND3X1_27 ( );
FILL FILL_1_NAND3X1_27 ( );
FILL FILL_2_NAND3X1_27 ( );
FILL FILL_3_NAND3X1_27 ( );
FILL FILL_4_NAND3X1_27 ( );
FILL FILL_5_NAND3X1_27 ( );
FILL FILL_6_NAND3X1_27 ( );
FILL FILL_7_NAND3X1_27 ( );
FILL FILL_8_NAND3X1_27 ( );
FILL FILL_9_NAND3X1_27 ( );
FILL FILL_0_NAND3X1_48 ( );
FILL FILL_1_NAND3X1_48 ( );
FILL FILL_2_NAND3X1_48 ( );
FILL FILL_3_NAND3X1_48 ( );
FILL FILL_4_NAND3X1_48 ( );
FILL FILL_5_NAND3X1_48 ( );
FILL FILL_6_NAND3X1_48 ( );
FILL FILL_7_NAND3X1_48 ( );
FILL FILL_8_NAND3X1_48 ( );
FILL FILL_9_NAND3X1_48 ( );
FILL FILL_0_NOR2X1_23 ( );
FILL FILL_1_NOR2X1_23 ( );
FILL FILL_2_NOR2X1_23 ( );
FILL FILL_3_NOR2X1_23 ( );
FILL FILL_4_NOR2X1_23 ( );
FILL FILL_5_NOR2X1_23 ( );
FILL FILL_6_NOR2X1_23 ( );
FILL FILL_0_NOR2X1_22 ( );
FILL FILL_1_NOR2X1_22 ( );
FILL FILL_2_NOR2X1_22 ( );
FILL FILL_3_NOR2X1_22 ( );
FILL FILL_4_NOR2X1_22 ( );
FILL FILL_5_NOR2X1_22 ( );
FILL FILL_6_NOR2X1_22 ( );
FILL FILL_0_CLKBUF1_9 ( );
FILL FILL_1_CLKBUF1_9 ( );
FILL FILL_2_CLKBUF1_9 ( );
FILL FILL_3_CLKBUF1_9 ( );
FILL FILL_4_CLKBUF1_9 ( );
FILL FILL_5_CLKBUF1_9 ( );
FILL FILL_6_CLKBUF1_9 ( );
FILL FILL_7_CLKBUF1_9 ( );
FILL FILL_8_CLKBUF1_9 ( );
FILL FILL_9_CLKBUF1_9 ( );
FILL FILL_10_CLKBUF1_9 ( );
FILL FILL_11_CLKBUF1_9 ( );
FILL FILL_12_CLKBUF1_9 ( );
FILL FILL_13_CLKBUF1_9 ( );
FILL FILL_14_CLKBUF1_9 ( );
FILL FILL_15_CLKBUF1_9 ( );
FILL FILL_16_CLKBUF1_9 ( );
FILL FILL_17_CLKBUF1_9 ( );
FILL FILL_18_CLKBUF1_9 ( );
FILL FILL_19_CLKBUF1_9 ( );
FILL FILL_20_CLKBUF1_9 ( );
FILL FILL_21_CLKBUF1_9 ( );
FILL FILL_0_DFFSR_119 ( );
FILL FILL_1_DFFSR_119 ( );
FILL FILL_2_DFFSR_119 ( );
FILL FILL_3_DFFSR_119 ( );
FILL FILL_4_DFFSR_119 ( );
FILL FILL_5_DFFSR_119 ( );
FILL FILL_6_DFFSR_119 ( );
FILL FILL_7_DFFSR_119 ( );
FILL FILL_8_DFFSR_119 ( );
FILL FILL_9_DFFSR_119 ( );
FILL FILL_10_DFFSR_119 ( );
FILL FILL_11_DFFSR_119 ( );
FILL FILL_12_DFFSR_119 ( );
FILL FILL_13_DFFSR_119 ( );
FILL FILL_14_DFFSR_119 ( );
FILL FILL_15_DFFSR_119 ( );
FILL FILL_16_DFFSR_119 ( );
FILL FILL_17_DFFSR_119 ( );
FILL FILL_18_DFFSR_119 ( );
FILL FILL_19_DFFSR_119 ( );
FILL FILL_20_DFFSR_119 ( );
FILL FILL_21_DFFSR_119 ( );
FILL FILL_22_DFFSR_119 ( );
FILL FILL_23_DFFSR_119 ( );
FILL FILL_24_DFFSR_119 ( );
FILL FILL_25_DFFSR_119 ( );
FILL FILL_26_DFFSR_119 ( );
FILL FILL_27_DFFSR_119 ( );
FILL FILL_28_DFFSR_119 ( );
FILL FILL_29_DFFSR_119 ( );
FILL FILL_30_DFFSR_119 ( );
FILL FILL_31_DFFSR_119 ( );
FILL FILL_32_DFFSR_119 ( );
FILL FILL_33_DFFSR_119 ( );
FILL FILL_34_DFFSR_119 ( );
FILL FILL_35_DFFSR_119 ( );
FILL FILL_36_DFFSR_119 ( );
FILL FILL_37_DFFSR_119 ( );
FILL FILL_38_DFFSR_119 ( );
FILL FILL_39_DFFSR_119 ( );
FILL FILL_40_DFFSR_119 ( );
FILL FILL_41_DFFSR_119 ( );
FILL FILL_42_DFFSR_119 ( );
FILL FILL_43_DFFSR_119 ( );
FILL FILL_44_DFFSR_119 ( );
FILL FILL_45_DFFSR_119 ( );
FILL FILL_46_DFFSR_119 ( );
FILL FILL_47_DFFSR_119 ( );
FILL FILL_48_DFFSR_119 ( );
FILL FILL_49_DFFSR_119 ( );
FILL FILL_50_DFFSR_119 ( );
FILL FILL_0_NOR2X1_18 ( );
FILL FILL_1_NOR2X1_18 ( );
FILL FILL_2_NOR2X1_18 ( );
FILL FILL_3_NOR2X1_18 ( );
FILL FILL_4_NOR2X1_18 ( );
FILL FILL_5_NOR2X1_18 ( );
FILL FILL_6_NOR2X1_18 ( );
FILL FILL_0_OAI22X1_14 ( );
FILL FILL_1_OAI22X1_14 ( );
FILL FILL_2_OAI22X1_14 ( );
FILL FILL_3_OAI22X1_14 ( );
FILL FILL_4_OAI22X1_14 ( );
FILL FILL_5_OAI22X1_14 ( );
FILL FILL_6_OAI22X1_14 ( );
FILL FILL_7_OAI22X1_14 ( );
FILL FILL_8_OAI22X1_14 ( );
FILL FILL_9_OAI22X1_14 ( );
FILL FILL_10_OAI22X1_14 ( );
FILL FILL_0_NAND3X1_40 ( );
FILL FILL_1_NAND3X1_40 ( );
FILL FILL_2_NAND3X1_40 ( );
FILL FILL_3_NAND3X1_40 ( );
FILL FILL_4_NAND3X1_40 ( );
FILL FILL_5_NAND3X1_40 ( );
FILL FILL_6_NAND3X1_40 ( );
FILL FILL_7_NAND3X1_40 ( );
FILL FILL_8_NAND3X1_40 ( );
FILL FILL_0_OAI21X1_6 ( );
FILL FILL_1_OAI21X1_6 ( );
FILL FILL_2_OAI21X1_6 ( );
FILL FILL_3_OAI21X1_6 ( );
FILL FILL_4_OAI21X1_6 ( );
FILL FILL_5_OAI21X1_6 ( );
FILL FILL_6_OAI21X1_6 ( );
FILL FILL_7_OAI21X1_6 ( );
FILL FILL_8_OAI21X1_6 ( );
FILL FILL_0_INVX1_44 ( );
FILL FILL_1_INVX1_44 ( );
FILL FILL_2_INVX1_44 ( );
FILL FILL_3_INVX1_44 ( );
FILL FILL_4_INVX1_44 ( );
FILL FILL_0_OAI22X1_9 ( );
FILL FILL_1_OAI22X1_9 ( );
FILL FILL_2_OAI22X1_9 ( );
FILL FILL_3_OAI22X1_9 ( );
FILL FILL_4_OAI22X1_9 ( );
FILL FILL_5_OAI22X1_9 ( );
FILL FILL_6_OAI22X1_9 ( );
FILL FILL_7_OAI22X1_9 ( );
FILL FILL_8_OAI22X1_9 ( );
FILL FILL_9_OAI22X1_9 ( );
FILL FILL_10_OAI22X1_9 ( );
FILL FILL_11_OAI22X1_9 ( );
FILL FILL_0_INVX1_34 ( );
FILL FILL_1_INVX1_34 ( );
FILL FILL_2_INVX1_34 ( );
FILL FILL_3_INVX1_34 ( );
FILL FILL_4_INVX1_34 ( );
FILL FILL_0_OAI22X1_3 ( );
FILL FILL_1_OAI22X1_3 ( );
FILL FILL_2_OAI22X1_3 ( );
FILL FILL_3_OAI22X1_3 ( );
FILL FILL_4_OAI22X1_3 ( );
FILL FILL_5_OAI22X1_3 ( );
FILL FILL_6_OAI22X1_3 ( );
FILL FILL_7_OAI22X1_3 ( );
FILL FILL_8_OAI22X1_3 ( );
FILL FILL_9_OAI22X1_3 ( );
FILL FILL_10_OAI22X1_3 ( );
FILL FILL_0_BUFX2_42 ( );
FILL FILL_1_BUFX2_42 ( );
FILL FILL_2_BUFX2_42 ( );
FILL FILL_3_BUFX2_42 ( );
FILL FILL_4_BUFX2_42 ( );
FILL FILL_5_BUFX2_42 ( );
FILL FILL_6_BUFX2_42 ( );
FILL FILL_0_INVX1_8 ( );
FILL FILL_1_INVX1_8 ( );
FILL FILL_2_INVX1_8 ( );
FILL FILL_3_INVX1_8 ( );
FILL FILL_4_INVX1_8 ( );
FILL FILL_0_DFFSR_25 ( );
FILL FILL_1_DFFSR_25 ( );
FILL FILL_2_DFFSR_25 ( );
FILL FILL_3_DFFSR_25 ( );
FILL FILL_4_DFFSR_25 ( );
FILL FILL_5_DFFSR_25 ( );
FILL FILL_6_DFFSR_25 ( );
FILL FILL_7_DFFSR_25 ( );
FILL FILL_8_DFFSR_25 ( );
FILL FILL_9_DFFSR_25 ( );
FILL FILL_10_DFFSR_25 ( );
FILL FILL_11_DFFSR_25 ( );
FILL FILL_12_DFFSR_25 ( );
FILL FILL_13_DFFSR_25 ( );
FILL FILL_14_DFFSR_25 ( );
FILL FILL_15_DFFSR_25 ( );
FILL FILL_16_DFFSR_25 ( );
FILL FILL_17_DFFSR_25 ( );
FILL FILL_18_DFFSR_25 ( );
FILL FILL_19_DFFSR_25 ( );
FILL FILL_20_DFFSR_25 ( );
FILL FILL_21_DFFSR_25 ( );
FILL FILL_22_DFFSR_25 ( );
FILL FILL_23_DFFSR_25 ( );
FILL FILL_24_DFFSR_25 ( );
FILL FILL_25_DFFSR_25 ( );
FILL FILL_26_DFFSR_25 ( );
FILL FILL_27_DFFSR_25 ( );
FILL FILL_28_DFFSR_25 ( );
FILL FILL_29_DFFSR_25 ( );
FILL FILL_30_DFFSR_25 ( );
FILL FILL_31_DFFSR_25 ( );
FILL FILL_32_DFFSR_25 ( );
FILL FILL_33_DFFSR_25 ( );
FILL FILL_34_DFFSR_25 ( );
FILL FILL_35_DFFSR_25 ( );
FILL FILL_36_DFFSR_25 ( );
FILL FILL_37_DFFSR_25 ( );
FILL FILL_38_DFFSR_25 ( );
FILL FILL_39_DFFSR_25 ( );
FILL FILL_40_DFFSR_25 ( );
FILL FILL_41_DFFSR_25 ( );
FILL FILL_42_DFFSR_25 ( );
FILL FILL_43_DFFSR_25 ( );
FILL FILL_44_DFFSR_25 ( );
FILL FILL_45_DFFSR_25 ( );
FILL FILL_46_DFFSR_25 ( );
FILL FILL_47_DFFSR_25 ( );
FILL FILL_48_DFFSR_25 ( );
FILL FILL_49_DFFSR_25 ( );
FILL FILL_50_DFFSR_25 ( );
FILL FILL_0_DFFSR_3 ( );
FILL FILL_1_DFFSR_3 ( );
FILL FILL_2_DFFSR_3 ( );
FILL FILL_3_DFFSR_3 ( );
FILL FILL_4_DFFSR_3 ( );
FILL FILL_5_DFFSR_3 ( );
FILL FILL_6_DFFSR_3 ( );
FILL FILL_7_DFFSR_3 ( );
FILL FILL_8_DFFSR_3 ( );
FILL FILL_9_DFFSR_3 ( );
FILL FILL_10_DFFSR_3 ( );
FILL FILL_11_DFFSR_3 ( );
FILL FILL_12_DFFSR_3 ( );
FILL FILL_13_DFFSR_3 ( );
FILL FILL_14_DFFSR_3 ( );
FILL FILL_15_DFFSR_3 ( );
FILL FILL_16_DFFSR_3 ( );
FILL FILL_17_DFFSR_3 ( );
FILL FILL_18_DFFSR_3 ( );
FILL FILL_19_DFFSR_3 ( );
FILL FILL_20_DFFSR_3 ( );
FILL FILL_21_DFFSR_3 ( );
FILL FILL_22_DFFSR_3 ( );
FILL FILL_23_DFFSR_3 ( );
FILL FILL_24_DFFSR_3 ( );
FILL FILL_25_DFFSR_3 ( );
FILL FILL_26_DFFSR_3 ( );
FILL FILL_27_DFFSR_3 ( );
FILL FILL_28_DFFSR_3 ( );
FILL FILL_29_DFFSR_3 ( );
FILL FILL_30_DFFSR_3 ( );
FILL FILL_31_DFFSR_3 ( );
FILL FILL_32_DFFSR_3 ( );
FILL FILL_33_DFFSR_3 ( );
FILL FILL_34_DFFSR_3 ( );
FILL FILL_35_DFFSR_3 ( );
FILL FILL_36_DFFSR_3 ( );
FILL FILL_37_DFFSR_3 ( );
FILL FILL_38_DFFSR_3 ( );
FILL FILL_39_DFFSR_3 ( );
FILL FILL_40_DFFSR_3 ( );
FILL FILL_41_DFFSR_3 ( );
FILL FILL_42_DFFSR_3 ( );
FILL FILL_43_DFFSR_3 ( );
FILL FILL_44_DFFSR_3 ( );
FILL FILL_45_DFFSR_3 ( );
FILL FILL_46_DFFSR_3 ( );
FILL FILL_47_DFFSR_3 ( );
FILL FILL_48_DFFSR_3 ( );
FILL FILL_49_DFFSR_3 ( );
FILL FILL_50_DFFSR_3 ( );
FILL FILL_51_DFFSR_3 ( );
FILL FILL_0_NAND3X1_242 ( );
FILL FILL_1_NAND3X1_242 ( );
FILL FILL_2_NAND3X1_242 ( );
FILL FILL_3_NAND3X1_242 ( );
FILL FILL_4_NAND3X1_242 ( );
FILL FILL_5_NAND3X1_242 ( );
FILL FILL_6_NAND3X1_242 ( );
FILL FILL_7_NAND3X1_242 ( );
FILL FILL_8_NAND3X1_242 ( );
FILL FILL_0_NAND3X1_243 ( );
FILL FILL_1_NAND3X1_243 ( );
FILL FILL_2_NAND3X1_243 ( );
FILL FILL_3_NAND3X1_243 ( );
FILL FILL_4_NAND3X1_243 ( );
FILL FILL_5_NAND3X1_243 ( );
FILL FILL_6_NAND3X1_243 ( );
FILL FILL_7_NAND3X1_243 ( );
FILL FILL_8_NAND3X1_243 ( );
FILL FILL_0_AOI21X1_44 ( );
FILL FILL_1_AOI21X1_44 ( );
FILL FILL_2_AOI21X1_44 ( );
FILL FILL_3_AOI21X1_44 ( );
FILL FILL_4_AOI21X1_44 ( );
FILL FILL_5_AOI21X1_44 ( );
FILL FILL_6_AOI21X1_44 ( );
FILL FILL_7_AOI21X1_44 ( );
FILL FILL_8_AOI21X1_44 ( );
FILL FILL_9_AOI21X1_44 ( );
FILL FILL_0_AOI21X1_45 ( );
FILL FILL_1_AOI21X1_45 ( );
FILL FILL_2_AOI21X1_45 ( );
FILL FILL_3_AOI21X1_45 ( );
FILL FILL_4_AOI21X1_45 ( );
FILL FILL_5_AOI21X1_45 ( );
FILL FILL_6_AOI21X1_45 ( );
FILL FILL_7_AOI21X1_45 ( );
FILL FILL_8_AOI21X1_45 ( );
FILL FILL_0_OAI22X1_52 ( );
FILL FILL_1_OAI22X1_52 ( );
FILL FILL_2_OAI22X1_52 ( );
FILL FILL_3_OAI22X1_52 ( );
FILL FILL_4_OAI22X1_52 ( );
FILL FILL_5_OAI22X1_52 ( );
FILL FILL_6_OAI22X1_52 ( );
FILL FILL_7_OAI22X1_52 ( );
FILL FILL_8_OAI22X1_52 ( );
FILL FILL_9_OAI22X1_52 ( );
FILL FILL_10_OAI22X1_52 ( );
FILL FILL_0_NAND2X1_115 ( );
FILL FILL_1_NAND2X1_115 ( );
FILL FILL_2_NAND2X1_115 ( );
FILL FILL_3_NAND2X1_115 ( );
FILL FILL_4_NAND2X1_115 ( );
FILL FILL_5_NAND2X1_115 ( );
FILL FILL_6_NAND2X1_115 ( );
FILL FILL_0_CLKBUF1_13 ( );
FILL FILL_1_CLKBUF1_13 ( );
FILL FILL_2_CLKBUF1_13 ( );
FILL FILL_3_CLKBUF1_13 ( );
FILL FILL_4_CLKBUF1_13 ( );
FILL FILL_5_CLKBUF1_13 ( );
FILL FILL_6_CLKBUF1_13 ( );
FILL FILL_7_CLKBUF1_13 ( );
FILL FILL_8_CLKBUF1_13 ( );
FILL FILL_9_CLKBUF1_13 ( );
FILL FILL_10_CLKBUF1_13 ( );
FILL FILL_11_CLKBUF1_13 ( );
FILL FILL_12_CLKBUF1_13 ( );
FILL FILL_13_CLKBUF1_13 ( );
FILL FILL_14_CLKBUF1_13 ( );
FILL FILL_15_CLKBUF1_13 ( );
FILL FILL_16_CLKBUF1_13 ( );
FILL FILL_17_CLKBUF1_13 ( );
FILL FILL_18_CLKBUF1_13 ( );
FILL FILL_19_CLKBUF1_13 ( );
FILL FILL_20_CLKBUF1_13 ( );
FILL FILL_0_DFFSR_58 ( );
FILL FILL_1_DFFSR_58 ( );
FILL FILL_2_DFFSR_58 ( );
FILL FILL_3_DFFSR_58 ( );
FILL FILL_4_DFFSR_58 ( );
FILL FILL_5_DFFSR_58 ( );
FILL FILL_6_DFFSR_58 ( );
FILL FILL_7_DFFSR_58 ( );
FILL FILL_8_DFFSR_58 ( );
FILL FILL_9_DFFSR_58 ( );
FILL FILL_10_DFFSR_58 ( );
FILL FILL_11_DFFSR_58 ( );
FILL FILL_12_DFFSR_58 ( );
FILL FILL_13_DFFSR_58 ( );
FILL FILL_14_DFFSR_58 ( );
FILL FILL_15_DFFSR_58 ( );
FILL FILL_16_DFFSR_58 ( );
FILL FILL_17_DFFSR_58 ( );
FILL FILL_18_DFFSR_58 ( );
FILL FILL_19_DFFSR_58 ( );
FILL FILL_20_DFFSR_58 ( );
FILL FILL_21_DFFSR_58 ( );
FILL FILL_22_DFFSR_58 ( );
FILL FILL_23_DFFSR_58 ( );
FILL FILL_24_DFFSR_58 ( );
FILL FILL_25_DFFSR_58 ( );
FILL FILL_26_DFFSR_58 ( );
FILL FILL_27_DFFSR_58 ( );
FILL FILL_28_DFFSR_58 ( );
FILL FILL_29_DFFSR_58 ( );
FILL FILL_30_DFFSR_58 ( );
FILL FILL_31_DFFSR_58 ( );
FILL FILL_32_DFFSR_58 ( );
FILL FILL_33_DFFSR_58 ( );
FILL FILL_34_DFFSR_58 ( );
FILL FILL_35_DFFSR_58 ( );
FILL FILL_36_DFFSR_58 ( );
FILL FILL_37_DFFSR_58 ( );
FILL FILL_38_DFFSR_58 ( );
FILL FILL_39_DFFSR_58 ( );
FILL FILL_40_DFFSR_58 ( );
FILL FILL_41_DFFSR_58 ( );
FILL FILL_42_DFFSR_58 ( );
FILL FILL_43_DFFSR_58 ( );
FILL FILL_44_DFFSR_58 ( );
FILL FILL_45_DFFSR_58 ( );
FILL FILL_46_DFFSR_58 ( );
FILL FILL_47_DFFSR_58 ( );
FILL FILL_48_DFFSR_58 ( );
FILL FILL_49_DFFSR_58 ( );
FILL FILL_50_DFFSR_58 ( );
FILL FILL_0_INVX1_28 ( );
FILL FILL_1_INVX1_28 ( );
FILL FILL_2_INVX1_28 ( );
FILL FILL_3_INVX1_28 ( );
FILL FILL_0_OAI22X1_12 ( );
FILL FILL_1_OAI22X1_12 ( );
FILL FILL_2_OAI22X1_12 ( );
FILL FILL_3_OAI22X1_12 ( );
FILL FILL_4_OAI22X1_12 ( );
FILL FILL_5_OAI22X1_12 ( );
FILL FILL_6_OAI22X1_12 ( );
FILL FILL_7_OAI22X1_12 ( );
FILL FILL_8_OAI22X1_12 ( );
FILL FILL_9_OAI22X1_12 ( );
FILL FILL_10_OAI22X1_12 ( );
FILL FILL_11_OAI22X1_12 ( );
FILL FILL_0_NAND3X1_58 ( );
FILL FILL_1_NAND3X1_58 ( );
FILL FILL_2_NAND3X1_58 ( );
FILL FILL_3_NAND3X1_58 ( );
FILL FILL_4_NAND3X1_58 ( );
FILL FILL_5_NAND3X1_58 ( );
FILL FILL_6_NAND3X1_58 ( );
FILL FILL_7_NAND3X1_58 ( );
FILL FILL_8_NAND3X1_58 ( );
FILL FILL_0_NAND3X1_26 ( );
FILL FILL_1_NAND3X1_26 ( );
FILL FILL_2_NAND3X1_26 ( );
FILL FILL_3_NAND3X1_26 ( );
FILL FILL_4_NAND3X1_26 ( );
FILL FILL_5_NAND3X1_26 ( );
FILL FILL_6_NAND3X1_26 ( );
FILL FILL_7_NAND3X1_26 ( );
FILL FILL_8_NAND3X1_26 ( );
FILL FILL_0_AND2X2_9 ( );
FILL FILL_1_AND2X2_9 ( );
FILL FILL_2_AND2X2_9 ( );
FILL FILL_3_AND2X2_9 ( );
FILL FILL_4_AND2X2_9 ( );
FILL FILL_5_AND2X2_9 ( );
FILL FILL_6_AND2X2_9 ( );
FILL FILL_7_AND2X2_9 ( );
FILL FILL_8_AND2X2_9 ( );
FILL FILL_0_NAND2X1_1 ( );
FILL FILL_1_NAND2X1_1 ( );
FILL FILL_2_NAND2X1_1 ( );
FILL FILL_3_NAND2X1_1 ( );
FILL FILL_4_NAND2X1_1 ( );
FILL FILL_5_NAND2X1_1 ( );
FILL FILL_6_NAND2X1_1 ( );
FILL FILL_0_AND2X2_13 ( );
FILL FILL_1_AND2X2_13 ( );
FILL FILL_2_AND2X2_13 ( );
FILL FILL_3_AND2X2_13 ( );
FILL FILL_4_AND2X2_13 ( );
FILL FILL_5_AND2X2_13 ( );
FILL FILL_6_AND2X2_13 ( );
FILL FILL_7_AND2X2_13 ( );
FILL FILL_8_AND2X2_13 ( );
FILL FILL_9_AND2X2_13 ( );
FILL FILL_0_BUFX2_19 ( );
FILL FILL_1_BUFX2_19 ( );
FILL FILL_2_BUFX2_19 ( );
FILL FILL_3_BUFX2_19 ( );
FILL FILL_4_BUFX2_19 ( );
FILL FILL_5_BUFX2_19 ( );
FILL FILL_6_BUFX2_19 ( );
FILL FILL_0_NOR2X1_21 ( );
FILL FILL_1_NOR2X1_21 ( );
FILL FILL_2_NOR2X1_21 ( );
FILL FILL_3_NOR2X1_21 ( );
FILL FILL_4_NOR2X1_21 ( );
FILL FILL_5_NOR2X1_21 ( );
FILL FILL_6_NOR2X1_21 ( );
FILL FILL_0_DFFSR_16 ( );
FILL FILL_1_DFFSR_16 ( );
FILL FILL_2_DFFSR_16 ( );
FILL FILL_3_DFFSR_16 ( );
FILL FILL_4_DFFSR_16 ( );
FILL FILL_5_DFFSR_16 ( );
FILL FILL_6_DFFSR_16 ( );
FILL FILL_7_DFFSR_16 ( );
FILL FILL_8_DFFSR_16 ( );
FILL FILL_9_DFFSR_16 ( );
FILL FILL_10_DFFSR_16 ( );
FILL FILL_11_DFFSR_16 ( );
FILL FILL_12_DFFSR_16 ( );
FILL FILL_13_DFFSR_16 ( );
FILL FILL_14_DFFSR_16 ( );
FILL FILL_15_DFFSR_16 ( );
FILL FILL_16_DFFSR_16 ( );
FILL FILL_17_DFFSR_16 ( );
FILL FILL_18_DFFSR_16 ( );
FILL FILL_19_DFFSR_16 ( );
FILL FILL_20_DFFSR_16 ( );
FILL FILL_21_DFFSR_16 ( );
FILL FILL_22_DFFSR_16 ( );
FILL FILL_23_DFFSR_16 ( );
FILL FILL_24_DFFSR_16 ( );
FILL FILL_25_DFFSR_16 ( );
FILL FILL_26_DFFSR_16 ( );
FILL FILL_27_DFFSR_16 ( );
FILL FILL_28_DFFSR_16 ( );
FILL FILL_29_DFFSR_16 ( );
FILL FILL_30_DFFSR_16 ( );
FILL FILL_31_DFFSR_16 ( );
FILL FILL_32_DFFSR_16 ( );
FILL FILL_33_DFFSR_16 ( );
FILL FILL_34_DFFSR_16 ( );
FILL FILL_35_DFFSR_16 ( );
FILL FILL_36_DFFSR_16 ( );
FILL FILL_37_DFFSR_16 ( );
FILL FILL_38_DFFSR_16 ( );
FILL FILL_39_DFFSR_16 ( );
FILL FILL_40_DFFSR_16 ( );
FILL FILL_41_DFFSR_16 ( );
FILL FILL_42_DFFSR_16 ( );
FILL FILL_43_DFFSR_16 ( );
FILL FILL_44_DFFSR_16 ( );
FILL FILL_45_DFFSR_16 ( );
FILL FILL_46_DFFSR_16 ( );
FILL FILL_47_DFFSR_16 ( );
FILL FILL_48_DFFSR_16 ( );
FILL FILL_49_DFFSR_16 ( );
FILL FILL_50_DFFSR_16 ( );
FILL FILL_0_NOR2X1_29 ( );
FILL FILL_1_NOR2X1_29 ( );
FILL FILL_2_NOR2X1_29 ( );
FILL FILL_3_NOR2X1_29 ( );
FILL FILL_4_NOR2X1_29 ( );
FILL FILL_5_NOR2X1_29 ( );
FILL FILL_6_NOR2X1_29 ( );
FILL FILL_0_NAND3X1_61 ( );
FILL FILL_1_NAND3X1_61 ( );
FILL FILL_2_NAND3X1_61 ( );
FILL FILL_3_NAND3X1_61 ( );
FILL FILL_4_NAND3X1_61 ( );
FILL FILL_5_NAND3X1_61 ( );
FILL FILL_6_NAND3X1_61 ( );
FILL FILL_7_NAND3X1_61 ( );
FILL FILL_8_NAND3X1_61 ( );
FILL FILL_0_NAND3X1_63 ( );
FILL FILL_1_NAND3X1_63 ( );
FILL FILL_2_NAND3X1_63 ( );
FILL FILL_3_NAND3X1_63 ( );
FILL FILL_4_NAND3X1_63 ( );
FILL FILL_5_NAND3X1_63 ( );
FILL FILL_6_NAND3X1_63 ( );
FILL FILL_7_NAND3X1_63 ( );
FILL FILL_8_NAND3X1_63 ( );
FILL FILL_9_NAND3X1_63 ( );
FILL FILL_0_DFFSR_35 ( );
FILL FILL_1_DFFSR_35 ( );
FILL FILL_2_DFFSR_35 ( );
FILL FILL_3_DFFSR_35 ( );
FILL FILL_4_DFFSR_35 ( );
FILL FILL_5_DFFSR_35 ( );
FILL FILL_6_DFFSR_35 ( );
FILL FILL_7_DFFSR_35 ( );
FILL FILL_8_DFFSR_35 ( );
FILL FILL_9_DFFSR_35 ( );
FILL FILL_10_DFFSR_35 ( );
FILL FILL_11_DFFSR_35 ( );
FILL FILL_12_DFFSR_35 ( );
FILL FILL_13_DFFSR_35 ( );
FILL FILL_14_DFFSR_35 ( );
FILL FILL_15_DFFSR_35 ( );
FILL FILL_16_DFFSR_35 ( );
FILL FILL_17_DFFSR_35 ( );
FILL FILL_18_DFFSR_35 ( );
FILL FILL_19_DFFSR_35 ( );
FILL FILL_20_DFFSR_35 ( );
FILL FILL_21_DFFSR_35 ( );
FILL FILL_22_DFFSR_35 ( );
FILL FILL_23_DFFSR_35 ( );
FILL FILL_24_DFFSR_35 ( );
FILL FILL_25_DFFSR_35 ( );
FILL FILL_26_DFFSR_35 ( );
FILL FILL_27_DFFSR_35 ( );
FILL FILL_28_DFFSR_35 ( );
FILL FILL_29_DFFSR_35 ( );
FILL FILL_30_DFFSR_35 ( );
FILL FILL_31_DFFSR_35 ( );
FILL FILL_32_DFFSR_35 ( );
FILL FILL_33_DFFSR_35 ( );
FILL FILL_34_DFFSR_35 ( );
FILL FILL_35_DFFSR_35 ( );
FILL FILL_36_DFFSR_35 ( );
FILL FILL_37_DFFSR_35 ( );
FILL FILL_38_DFFSR_35 ( );
FILL FILL_39_DFFSR_35 ( );
FILL FILL_40_DFFSR_35 ( );
FILL FILL_41_DFFSR_35 ( );
FILL FILL_42_DFFSR_35 ( );
FILL FILL_43_DFFSR_35 ( );
FILL FILL_44_DFFSR_35 ( );
FILL FILL_45_DFFSR_35 ( );
FILL FILL_46_DFFSR_35 ( );
FILL FILL_47_DFFSR_35 ( );
FILL FILL_48_DFFSR_35 ( );
FILL FILL_49_DFFSR_35 ( );
FILL FILL_50_DFFSR_35 ( );
FILL FILL_0_INVX1_33 ( );
FILL FILL_1_INVX1_33 ( );
FILL FILL_2_INVX1_33 ( );
FILL FILL_3_INVX1_33 ( );
FILL FILL_4_INVX1_33 ( );
FILL FILL_0_NOR2X1_19 ( );
FILL FILL_1_NOR2X1_19 ( );
FILL FILL_2_NOR2X1_19 ( );
FILL FILL_3_NOR2X1_19 ( );
FILL FILL_4_NOR2X1_19 ( );
FILL FILL_5_NOR2X1_19 ( );
FILL FILL_6_NOR2X1_19 ( );
FILL FILL_0_OAI22X1_15 ( );
FILL FILL_1_OAI22X1_15 ( );
FILL FILL_2_OAI22X1_15 ( );
FILL FILL_3_OAI22X1_15 ( );
FILL FILL_4_OAI22X1_15 ( );
FILL FILL_5_OAI22X1_15 ( );
FILL FILL_6_OAI22X1_15 ( );
FILL FILL_7_OAI22X1_15 ( );
FILL FILL_8_OAI22X1_15 ( );
FILL FILL_9_OAI22X1_15 ( );
FILL FILL_10_OAI22X1_15 ( );
FILL FILL_0_INVX1_35 ( );
FILL FILL_1_INVX1_35 ( );
FILL FILL_2_INVX1_35 ( );
FILL FILL_3_INVX1_35 ( );
FILL FILL_4_INVX1_35 ( );
FILL FILL_0_AOI22X1_8 ( );
FILL FILL_1_AOI22X1_8 ( );
FILL FILL_2_AOI22X1_8 ( );
FILL FILL_3_AOI22X1_8 ( );
FILL FILL_4_AOI22X1_8 ( );
FILL FILL_5_AOI22X1_8 ( );
FILL FILL_6_AOI22X1_8 ( );
FILL FILL_7_AOI22X1_8 ( );
FILL FILL_8_AOI22X1_8 ( );
FILL FILL_9_AOI22X1_8 ( );
FILL FILL_10_AOI22X1_8 ( );
FILL FILL_0_DFFSR_17 ( );
FILL FILL_1_DFFSR_17 ( );
FILL FILL_2_DFFSR_17 ( );
FILL FILL_3_DFFSR_17 ( );
FILL FILL_4_DFFSR_17 ( );
FILL FILL_5_DFFSR_17 ( );
FILL FILL_6_DFFSR_17 ( );
FILL FILL_7_DFFSR_17 ( );
FILL FILL_8_DFFSR_17 ( );
FILL FILL_9_DFFSR_17 ( );
FILL FILL_10_DFFSR_17 ( );
FILL FILL_11_DFFSR_17 ( );
FILL FILL_12_DFFSR_17 ( );
FILL FILL_13_DFFSR_17 ( );
FILL FILL_14_DFFSR_17 ( );
FILL FILL_15_DFFSR_17 ( );
FILL FILL_16_DFFSR_17 ( );
FILL FILL_17_DFFSR_17 ( );
FILL FILL_18_DFFSR_17 ( );
FILL FILL_19_DFFSR_17 ( );
FILL FILL_20_DFFSR_17 ( );
FILL FILL_21_DFFSR_17 ( );
FILL FILL_22_DFFSR_17 ( );
FILL FILL_23_DFFSR_17 ( );
FILL FILL_24_DFFSR_17 ( );
FILL FILL_25_DFFSR_17 ( );
FILL FILL_26_DFFSR_17 ( );
FILL FILL_27_DFFSR_17 ( );
FILL FILL_28_DFFSR_17 ( );
FILL FILL_29_DFFSR_17 ( );
FILL FILL_30_DFFSR_17 ( );
FILL FILL_31_DFFSR_17 ( );
FILL FILL_32_DFFSR_17 ( );
FILL FILL_33_DFFSR_17 ( );
FILL FILL_34_DFFSR_17 ( );
FILL FILL_35_DFFSR_17 ( );
FILL FILL_36_DFFSR_17 ( );
FILL FILL_37_DFFSR_17 ( );
FILL FILL_38_DFFSR_17 ( );
FILL FILL_39_DFFSR_17 ( );
FILL FILL_40_DFFSR_17 ( );
FILL FILL_41_DFFSR_17 ( );
FILL FILL_42_DFFSR_17 ( );
FILL FILL_43_DFFSR_17 ( );
FILL FILL_44_DFFSR_17 ( );
FILL FILL_45_DFFSR_17 ( );
FILL FILL_46_DFFSR_17 ( );
FILL FILL_47_DFFSR_17 ( );
FILL FILL_48_DFFSR_17 ( );
FILL FILL_49_DFFSR_17 ( );
FILL FILL_50_DFFSR_17 ( );
FILL FILL_51_DFFSR_17 ( );
FILL FILL_0_BUFX2_91 ( );
FILL FILL_1_BUFX2_91 ( );
FILL FILL_2_BUFX2_91 ( );
FILL FILL_3_BUFX2_91 ( );
FILL FILL_4_BUFX2_91 ( );
FILL FILL_5_BUFX2_91 ( );
FILL FILL_6_BUFX2_91 ( );
FILL FILL_0_DFFSR_27 ( );
FILL FILL_1_DFFSR_27 ( );
FILL FILL_2_DFFSR_27 ( );
FILL FILL_3_DFFSR_27 ( );
FILL FILL_4_DFFSR_27 ( );
FILL FILL_5_DFFSR_27 ( );
FILL FILL_6_DFFSR_27 ( );
FILL FILL_7_DFFSR_27 ( );
FILL FILL_8_DFFSR_27 ( );
FILL FILL_9_DFFSR_27 ( );
FILL FILL_10_DFFSR_27 ( );
FILL FILL_11_DFFSR_27 ( );
FILL FILL_12_DFFSR_27 ( );
FILL FILL_13_DFFSR_27 ( );
FILL FILL_14_DFFSR_27 ( );
FILL FILL_15_DFFSR_27 ( );
FILL FILL_16_DFFSR_27 ( );
FILL FILL_17_DFFSR_27 ( );
FILL FILL_18_DFFSR_27 ( );
FILL FILL_19_DFFSR_27 ( );
FILL FILL_20_DFFSR_27 ( );
FILL FILL_21_DFFSR_27 ( );
FILL FILL_22_DFFSR_27 ( );
FILL FILL_23_DFFSR_27 ( );
FILL FILL_24_DFFSR_27 ( );
FILL FILL_25_DFFSR_27 ( );
FILL FILL_26_DFFSR_27 ( );
FILL FILL_27_DFFSR_27 ( );
FILL FILL_28_DFFSR_27 ( );
FILL FILL_29_DFFSR_27 ( );
FILL FILL_30_DFFSR_27 ( );
FILL FILL_31_DFFSR_27 ( );
FILL FILL_32_DFFSR_27 ( );
FILL FILL_33_DFFSR_27 ( );
FILL FILL_34_DFFSR_27 ( );
FILL FILL_35_DFFSR_27 ( );
FILL FILL_36_DFFSR_27 ( );
FILL FILL_37_DFFSR_27 ( );
FILL FILL_38_DFFSR_27 ( );
FILL FILL_39_DFFSR_27 ( );
FILL FILL_40_DFFSR_27 ( );
FILL FILL_41_DFFSR_27 ( );
FILL FILL_42_DFFSR_27 ( );
FILL FILL_43_DFFSR_27 ( );
FILL FILL_44_DFFSR_27 ( );
FILL FILL_45_DFFSR_27 ( );
FILL FILL_46_DFFSR_27 ( );
FILL FILL_47_DFFSR_27 ( );
FILL FILL_48_DFFSR_27 ( );
FILL FILL_49_DFFSR_27 ( );
FILL FILL_50_DFFSR_27 ( );
FILL FILL_51_DFFSR_27 ( );
FILL FILL_0_INVX1_172 ( );
FILL FILL_1_INVX1_172 ( );
FILL FILL_2_INVX1_172 ( );
FILL FILL_3_INVX1_172 ( );
FILL FILL_4_INVX1_172 ( );
FILL FILL_0_AOI21X1_38 ( );
FILL FILL_1_AOI21X1_38 ( );
FILL FILL_2_AOI21X1_38 ( );
FILL FILL_3_AOI21X1_38 ( );
FILL FILL_4_AOI21X1_38 ( );
FILL FILL_5_AOI21X1_38 ( );
FILL FILL_6_AOI21X1_38 ( );
FILL FILL_7_AOI21X1_38 ( );
FILL FILL_8_AOI21X1_38 ( );
FILL FILL_0_OAI21X1_82 ( );
FILL FILL_1_OAI21X1_82 ( );
FILL FILL_2_OAI21X1_82 ( );
FILL FILL_3_OAI21X1_82 ( );
FILL FILL_4_OAI21X1_82 ( );
FILL FILL_5_OAI21X1_82 ( );
FILL FILL_6_OAI21X1_82 ( );
FILL FILL_7_OAI21X1_82 ( );
FILL FILL_8_OAI21X1_82 ( );
FILL FILL_0_INVX1_170 ( );
FILL FILL_1_INVX1_170 ( );
FILL FILL_2_INVX1_170 ( );
FILL FILL_3_INVX1_170 ( );
FILL FILL_0_NAND3X1_244 ( );
FILL FILL_1_NAND3X1_244 ( );
FILL FILL_2_NAND3X1_244 ( );
FILL FILL_3_NAND3X1_244 ( );
FILL FILL_4_NAND3X1_244 ( );
FILL FILL_5_NAND3X1_244 ( );
FILL FILL_6_NAND3X1_244 ( );
FILL FILL_7_NAND3X1_244 ( );
FILL FILL_8_NAND3X1_244 ( );
FILL FILL_9_NAND3X1_244 ( );
FILL FILL_0_DFFPOSX1_21 ( );
FILL FILL_1_DFFPOSX1_21 ( );
FILL FILL_2_DFFPOSX1_21 ( );
FILL FILL_3_DFFPOSX1_21 ( );
FILL FILL_4_DFFPOSX1_21 ( );
FILL FILL_5_DFFPOSX1_21 ( );
FILL FILL_6_DFFPOSX1_21 ( );
FILL FILL_7_DFFPOSX1_21 ( );
FILL FILL_8_DFFPOSX1_21 ( );
FILL FILL_9_DFFPOSX1_21 ( );
FILL FILL_10_DFFPOSX1_21 ( );
FILL FILL_11_DFFPOSX1_21 ( );
FILL FILL_12_DFFPOSX1_21 ( );
FILL FILL_13_DFFPOSX1_21 ( );
FILL FILL_14_DFFPOSX1_21 ( );
FILL FILL_15_DFFPOSX1_21 ( );
FILL FILL_16_DFFPOSX1_21 ( );
FILL FILL_17_DFFPOSX1_21 ( );
FILL FILL_18_DFFPOSX1_21 ( );
FILL FILL_19_DFFPOSX1_21 ( );
FILL FILL_20_DFFPOSX1_21 ( );
FILL FILL_21_DFFPOSX1_21 ( );
FILL FILL_22_DFFPOSX1_21 ( );
FILL FILL_23_DFFPOSX1_21 ( );
FILL FILL_24_DFFPOSX1_21 ( );
FILL FILL_25_DFFPOSX1_21 ( );
FILL FILL_26_DFFPOSX1_21 ( );
FILL FILL_27_DFFPOSX1_21 ( );
FILL FILL_0_DFFSR_28 ( );
FILL FILL_1_DFFSR_28 ( );
FILL FILL_2_DFFSR_28 ( );
FILL FILL_3_DFFSR_28 ( );
FILL FILL_4_DFFSR_28 ( );
FILL FILL_5_DFFSR_28 ( );
FILL FILL_6_DFFSR_28 ( );
FILL FILL_7_DFFSR_28 ( );
FILL FILL_8_DFFSR_28 ( );
FILL FILL_9_DFFSR_28 ( );
FILL FILL_10_DFFSR_28 ( );
FILL FILL_11_DFFSR_28 ( );
FILL FILL_12_DFFSR_28 ( );
FILL FILL_13_DFFSR_28 ( );
FILL FILL_14_DFFSR_28 ( );
FILL FILL_15_DFFSR_28 ( );
FILL FILL_16_DFFSR_28 ( );
FILL FILL_17_DFFSR_28 ( );
FILL FILL_18_DFFSR_28 ( );
FILL FILL_19_DFFSR_28 ( );
FILL FILL_20_DFFSR_28 ( );
FILL FILL_21_DFFSR_28 ( );
FILL FILL_22_DFFSR_28 ( );
FILL FILL_23_DFFSR_28 ( );
FILL FILL_24_DFFSR_28 ( );
FILL FILL_25_DFFSR_28 ( );
FILL FILL_26_DFFSR_28 ( );
FILL FILL_27_DFFSR_28 ( );
FILL FILL_28_DFFSR_28 ( );
FILL FILL_29_DFFSR_28 ( );
FILL FILL_30_DFFSR_28 ( );
FILL FILL_31_DFFSR_28 ( );
FILL FILL_32_DFFSR_28 ( );
FILL FILL_33_DFFSR_28 ( );
FILL FILL_34_DFFSR_28 ( );
FILL FILL_35_DFFSR_28 ( );
FILL FILL_36_DFFSR_28 ( );
FILL FILL_37_DFFSR_28 ( );
FILL FILL_38_DFFSR_28 ( );
FILL FILL_39_DFFSR_28 ( );
FILL FILL_40_DFFSR_28 ( );
FILL FILL_41_DFFSR_28 ( );
FILL FILL_42_DFFSR_28 ( );
FILL FILL_43_DFFSR_28 ( );
FILL FILL_44_DFFSR_28 ( );
FILL FILL_45_DFFSR_28 ( );
FILL FILL_46_DFFSR_28 ( );
FILL FILL_47_DFFSR_28 ( );
FILL FILL_48_DFFSR_28 ( );
FILL FILL_49_DFFSR_28 ( );
FILL FILL_50_DFFSR_28 ( );
FILL FILL_0_INVX1_29 ( );
FILL FILL_1_INVX1_29 ( );
FILL FILL_2_INVX1_29 ( );
FILL FILL_3_INVX1_29 ( );
FILL FILL_4_INVX1_29 ( );
FILL FILL_0_DFFSR_56 ( );
FILL FILL_1_DFFSR_56 ( );
FILL FILL_2_DFFSR_56 ( );
FILL FILL_3_DFFSR_56 ( );
FILL FILL_4_DFFSR_56 ( );
FILL FILL_5_DFFSR_56 ( );
FILL FILL_6_DFFSR_56 ( );
FILL FILL_7_DFFSR_56 ( );
FILL FILL_8_DFFSR_56 ( );
FILL FILL_9_DFFSR_56 ( );
FILL FILL_10_DFFSR_56 ( );
FILL FILL_11_DFFSR_56 ( );
FILL FILL_12_DFFSR_56 ( );
FILL FILL_13_DFFSR_56 ( );
FILL FILL_14_DFFSR_56 ( );
FILL FILL_15_DFFSR_56 ( );
FILL FILL_16_DFFSR_56 ( );
FILL FILL_17_DFFSR_56 ( );
FILL FILL_18_DFFSR_56 ( );
FILL FILL_19_DFFSR_56 ( );
FILL FILL_20_DFFSR_56 ( );
FILL FILL_21_DFFSR_56 ( );
FILL FILL_22_DFFSR_56 ( );
FILL FILL_23_DFFSR_56 ( );
FILL FILL_24_DFFSR_56 ( );
FILL FILL_25_DFFSR_56 ( );
FILL FILL_26_DFFSR_56 ( );
FILL FILL_27_DFFSR_56 ( );
FILL FILL_28_DFFSR_56 ( );
FILL FILL_29_DFFSR_56 ( );
FILL FILL_30_DFFSR_56 ( );
FILL FILL_31_DFFSR_56 ( );
FILL FILL_32_DFFSR_56 ( );
FILL FILL_33_DFFSR_56 ( );
FILL FILL_34_DFFSR_56 ( );
FILL FILL_35_DFFSR_56 ( );
FILL FILL_36_DFFSR_56 ( );
FILL FILL_37_DFFSR_56 ( );
FILL FILL_38_DFFSR_56 ( );
FILL FILL_39_DFFSR_56 ( );
FILL FILL_40_DFFSR_56 ( );
FILL FILL_41_DFFSR_56 ( );
FILL FILL_42_DFFSR_56 ( );
FILL FILL_43_DFFSR_56 ( );
FILL FILL_44_DFFSR_56 ( );
FILL FILL_45_DFFSR_56 ( );
FILL FILL_46_DFFSR_56 ( );
FILL FILL_47_DFFSR_56 ( );
FILL FILL_48_DFFSR_56 ( );
FILL FILL_49_DFFSR_56 ( );
FILL FILL_50_DFFSR_56 ( );
FILL FILL_0_BUFX2_12 ( );
FILL FILL_1_BUFX2_12 ( );
FILL FILL_2_BUFX2_12 ( );
FILL FILL_3_BUFX2_12 ( );
FILL FILL_4_BUFX2_12 ( );
FILL FILL_5_BUFX2_12 ( );
FILL FILL_6_BUFX2_12 ( );
FILL FILL_0_BUFX2_13 ( );
FILL FILL_1_BUFX2_13 ( );
FILL FILL_2_BUFX2_13 ( );
FILL FILL_3_BUFX2_13 ( );
FILL FILL_4_BUFX2_13 ( );
FILL FILL_5_BUFX2_13 ( );
FILL FILL_6_BUFX2_13 ( );
FILL FILL_0_NAND3X1_56 ( );
FILL FILL_1_NAND3X1_56 ( );
FILL FILL_2_NAND3X1_56 ( );
FILL FILL_3_NAND3X1_56 ( );
FILL FILL_4_NAND3X1_56 ( );
FILL FILL_5_NAND3X1_56 ( );
FILL FILL_6_NAND3X1_56 ( );
FILL FILL_7_NAND3X1_56 ( );
FILL FILL_8_NAND3X1_56 ( );
FILL FILL_0_NAND3X1_16 ( );
FILL FILL_1_NAND3X1_16 ( );
FILL FILL_2_NAND3X1_16 ( );
FILL FILL_3_NAND3X1_16 ( );
FILL FILL_4_NAND3X1_16 ( );
FILL FILL_5_NAND3X1_16 ( );
FILL FILL_6_NAND3X1_16 ( );
FILL FILL_7_NAND3X1_16 ( );
FILL FILL_8_NAND3X1_16 ( );
FILL FILL_0_NOR2X1_25 ( );
FILL FILL_1_NOR2X1_25 ( );
FILL FILL_2_NOR2X1_25 ( );
FILL FILL_3_NOR2X1_25 ( );
FILL FILL_4_NOR2X1_25 ( );
FILL FILL_5_NOR2X1_25 ( );
FILL FILL_6_NOR2X1_25 ( );
FILL FILL_0_INVX1_51 ( );
FILL FILL_1_INVX1_51 ( );
FILL FILL_2_INVX1_51 ( );
FILL FILL_3_INVX1_51 ( );
FILL FILL_0_DFFSR_70 ( );
FILL FILL_1_DFFSR_70 ( );
FILL FILL_2_DFFSR_70 ( );
FILL FILL_3_DFFSR_70 ( );
FILL FILL_4_DFFSR_70 ( );
FILL FILL_5_DFFSR_70 ( );
FILL FILL_6_DFFSR_70 ( );
FILL FILL_7_DFFSR_70 ( );
FILL FILL_8_DFFSR_70 ( );
FILL FILL_9_DFFSR_70 ( );
FILL FILL_10_DFFSR_70 ( );
FILL FILL_11_DFFSR_70 ( );
FILL FILL_12_DFFSR_70 ( );
FILL FILL_13_DFFSR_70 ( );
FILL FILL_14_DFFSR_70 ( );
FILL FILL_15_DFFSR_70 ( );
FILL FILL_16_DFFSR_70 ( );
FILL FILL_17_DFFSR_70 ( );
FILL FILL_18_DFFSR_70 ( );
FILL FILL_19_DFFSR_70 ( );
FILL FILL_20_DFFSR_70 ( );
FILL FILL_21_DFFSR_70 ( );
FILL FILL_22_DFFSR_70 ( );
FILL FILL_23_DFFSR_70 ( );
FILL FILL_24_DFFSR_70 ( );
FILL FILL_25_DFFSR_70 ( );
FILL FILL_26_DFFSR_70 ( );
FILL FILL_27_DFFSR_70 ( );
FILL FILL_28_DFFSR_70 ( );
FILL FILL_29_DFFSR_70 ( );
FILL FILL_30_DFFSR_70 ( );
FILL FILL_31_DFFSR_70 ( );
FILL FILL_32_DFFSR_70 ( );
FILL FILL_33_DFFSR_70 ( );
FILL FILL_34_DFFSR_70 ( );
FILL FILL_35_DFFSR_70 ( );
FILL FILL_36_DFFSR_70 ( );
FILL FILL_37_DFFSR_70 ( );
FILL FILL_38_DFFSR_70 ( );
FILL FILL_39_DFFSR_70 ( );
FILL FILL_40_DFFSR_70 ( );
FILL FILL_41_DFFSR_70 ( );
FILL FILL_42_DFFSR_70 ( );
FILL FILL_43_DFFSR_70 ( );
FILL FILL_44_DFFSR_70 ( );
FILL FILL_45_DFFSR_70 ( );
FILL FILL_46_DFFSR_70 ( );
FILL FILL_47_DFFSR_70 ( );
FILL FILL_48_DFFSR_70 ( );
FILL FILL_49_DFFSR_70 ( );
FILL FILL_50_DFFSR_70 ( );
FILL FILL_0_DFFSR_61 ( );
FILL FILL_1_DFFSR_61 ( );
FILL FILL_2_DFFSR_61 ( );
FILL FILL_3_DFFSR_61 ( );
FILL FILL_4_DFFSR_61 ( );
FILL FILL_5_DFFSR_61 ( );
FILL FILL_6_DFFSR_61 ( );
FILL FILL_7_DFFSR_61 ( );
FILL FILL_8_DFFSR_61 ( );
FILL FILL_9_DFFSR_61 ( );
FILL FILL_10_DFFSR_61 ( );
FILL FILL_11_DFFSR_61 ( );
FILL FILL_12_DFFSR_61 ( );
FILL FILL_13_DFFSR_61 ( );
FILL FILL_14_DFFSR_61 ( );
FILL FILL_15_DFFSR_61 ( );
FILL FILL_16_DFFSR_61 ( );
FILL FILL_17_DFFSR_61 ( );
FILL FILL_18_DFFSR_61 ( );
FILL FILL_19_DFFSR_61 ( );
FILL FILL_20_DFFSR_61 ( );
FILL FILL_21_DFFSR_61 ( );
FILL FILL_22_DFFSR_61 ( );
FILL FILL_23_DFFSR_61 ( );
FILL FILL_24_DFFSR_61 ( );
FILL FILL_25_DFFSR_61 ( );
FILL FILL_26_DFFSR_61 ( );
FILL FILL_27_DFFSR_61 ( );
FILL FILL_28_DFFSR_61 ( );
FILL FILL_29_DFFSR_61 ( );
FILL FILL_30_DFFSR_61 ( );
FILL FILL_31_DFFSR_61 ( );
FILL FILL_32_DFFSR_61 ( );
FILL FILL_33_DFFSR_61 ( );
FILL FILL_34_DFFSR_61 ( );
FILL FILL_35_DFFSR_61 ( );
FILL FILL_36_DFFSR_61 ( );
FILL FILL_37_DFFSR_61 ( );
FILL FILL_38_DFFSR_61 ( );
FILL FILL_39_DFFSR_61 ( );
FILL FILL_40_DFFSR_61 ( );
FILL FILL_41_DFFSR_61 ( );
FILL FILL_42_DFFSR_61 ( );
FILL FILL_43_DFFSR_61 ( );
FILL FILL_44_DFFSR_61 ( );
FILL FILL_45_DFFSR_61 ( );
FILL FILL_46_DFFSR_61 ( );
FILL FILL_47_DFFSR_61 ( );
FILL FILL_48_DFFSR_61 ( );
FILL FILL_49_DFFSR_61 ( );
FILL FILL_50_DFFSR_61 ( );
FILL FILL_0_NAND2X1_21 ( );
FILL FILL_1_NAND2X1_21 ( );
FILL FILL_2_NAND2X1_21 ( );
FILL FILL_3_NAND2X1_21 ( );
FILL FILL_4_NAND2X1_21 ( );
FILL FILL_5_NAND2X1_21 ( );
FILL FILL_6_NAND2X1_21 ( );
FILL FILL_0_DFFSR_104 ( );
FILL FILL_1_DFFSR_104 ( );
FILL FILL_2_DFFSR_104 ( );
FILL FILL_3_DFFSR_104 ( );
FILL FILL_4_DFFSR_104 ( );
FILL FILL_5_DFFSR_104 ( );
FILL FILL_6_DFFSR_104 ( );
FILL FILL_7_DFFSR_104 ( );
FILL FILL_8_DFFSR_104 ( );
FILL FILL_9_DFFSR_104 ( );
FILL FILL_10_DFFSR_104 ( );
FILL FILL_11_DFFSR_104 ( );
FILL FILL_12_DFFSR_104 ( );
FILL FILL_13_DFFSR_104 ( );
FILL FILL_14_DFFSR_104 ( );
FILL FILL_15_DFFSR_104 ( );
FILL FILL_16_DFFSR_104 ( );
FILL FILL_17_DFFSR_104 ( );
FILL FILL_18_DFFSR_104 ( );
FILL FILL_19_DFFSR_104 ( );
FILL FILL_20_DFFSR_104 ( );
FILL FILL_21_DFFSR_104 ( );
FILL FILL_22_DFFSR_104 ( );
FILL FILL_23_DFFSR_104 ( );
FILL FILL_24_DFFSR_104 ( );
FILL FILL_25_DFFSR_104 ( );
FILL FILL_26_DFFSR_104 ( );
FILL FILL_27_DFFSR_104 ( );
FILL FILL_28_DFFSR_104 ( );
FILL FILL_29_DFFSR_104 ( );
FILL FILL_30_DFFSR_104 ( );
FILL FILL_31_DFFSR_104 ( );
FILL FILL_32_DFFSR_104 ( );
FILL FILL_33_DFFSR_104 ( );
FILL FILL_34_DFFSR_104 ( );
FILL FILL_35_DFFSR_104 ( );
FILL FILL_36_DFFSR_104 ( );
FILL FILL_37_DFFSR_104 ( );
FILL FILL_38_DFFSR_104 ( );
FILL FILL_39_DFFSR_104 ( );
FILL FILL_40_DFFSR_104 ( );
FILL FILL_41_DFFSR_104 ( );
FILL FILL_42_DFFSR_104 ( );
FILL FILL_43_DFFSR_104 ( );
FILL FILL_44_DFFSR_104 ( );
FILL FILL_45_DFFSR_104 ( );
FILL FILL_46_DFFSR_104 ( );
FILL FILL_47_DFFSR_104 ( );
FILL FILL_48_DFFSR_104 ( );
FILL FILL_49_DFFSR_104 ( );
FILL FILL_50_DFFSR_104 ( );
FILL FILL_0_DFFSR_19 ( );
FILL FILL_1_DFFSR_19 ( );
FILL FILL_2_DFFSR_19 ( );
FILL FILL_3_DFFSR_19 ( );
FILL FILL_4_DFFSR_19 ( );
FILL FILL_5_DFFSR_19 ( );
FILL FILL_6_DFFSR_19 ( );
FILL FILL_7_DFFSR_19 ( );
FILL FILL_8_DFFSR_19 ( );
FILL FILL_9_DFFSR_19 ( );
FILL FILL_10_DFFSR_19 ( );
FILL FILL_11_DFFSR_19 ( );
FILL FILL_12_DFFSR_19 ( );
FILL FILL_13_DFFSR_19 ( );
FILL FILL_14_DFFSR_19 ( );
FILL FILL_15_DFFSR_19 ( );
FILL FILL_16_DFFSR_19 ( );
FILL FILL_17_DFFSR_19 ( );
FILL FILL_18_DFFSR_19 ( );
FILL FILL_19_DFFSR_19 ( );
FILL FILL_20_DFFSR_19 ( );
FILL FILL_21_DFFSR_19 ( );
FILL FILL_22_DFFSR_19 ( );
FILL FILL_23_DFFSR_19 ( );
FILL FILL_24_DFFSR_19 ( );
FILL FILL_25_DFFSR_19 ( );
FILL FILL_26_DFFSR_19 ( );
FILL FILL_27_DFFSR_19 ( );
FILL FILL_28_DFFSR_19 ( );
FILL FILL_29_DFFSR_19 ( );
FILL FILL_30_DFFSR_19 ( );
FILL FILL_31_DFFSR_19 ( );
FILL FILL_32_DFFSR_19 ( );
FILL FILL_33_DFFSR_19 ( );
FILL FILL_34_DFFSR_19 ( );
FILL FILL_35_DFFSR_19 ( );
FILL FILL_36_DFFSR_19 ( );
FILL FILL_37_DFFSR_19 ( );
FILL FILL_38_DFFSR_19 ( );
FILL FILL_39_DFFSR_19 ( );
FILL FILL_40_DFFSR_19 ( );
FILL FILL_41_DFFSR_19 ( );
FILL FILL_42_DFFSR_19 ( );
FILL FILL_43_DFFSR_19 ( );
FILL FILL_44_DFFSR_19 ( );
FILL FILL_45_DFFSR_19 ( );
FILL FILL_46_DFFSR_19 ( );
FILL FILL_47_DFFSR_19 ( );
FILL FILL_48_DFFSR_19 ( );
FILL FILL_49_DFFSR_19 ( );
FILL FILL_50_DFFSR_19 ( );
FILL FILL_0_DFFSR_248 ( );
FILL FILL_1_DFFSR_248 ( );
FILL FILL_2_DFFSR_248 ( );
FILL FILL_3_DFFSR_248 ( );
FILL FILL_4_DFFSR_248 ( );
FILL FILL_5_DFFSR_248 ( );
FILL FILL_6_DFFSR_248 ( );
FILL FILL_7_DFFSR_248 ( );
FILL FILL_8_DFFSR_248 ( );
FILL FILL_9_DFFSR_248 ( );
FILL FILL_10_DFFSR_248 ( );
FILL FILL_11_DFFSR_248 ( );
FILL FILL_12_DFFSR_248 ( );
FILL FILL_13_DFFSR_248 ( );
FILL FILL_14_DFFSR_248 ( );
FILL FILL_15_DFFSR_248 ( );
FILL FILL_16_DFFSR_248 ( );
FILL FILL_17_DFFSR_248 ( );
FILL FILL_18_DFFSR_248 ( );
FILL FILL_19_DFFSR_248 ( );
FILL FILL_20_DFFSR_248 ( );
FILL FILL_21_DFFSR_248 ( );
FILL FILL_22_DFFSR_248 ( );
FILL FILL_23_DFFSR_248 ( );
FILL FILL_24_DFFSR_248 ( );
FILL FILL_25_DFFSR_248 ( );
FILL FILL_26_DFFSR_248 ( );
FILL FILL_27_DFFSR_248 ( );
FILL FILL_28_DFFSR_248 ( );
FILL FILL_29_DFFSR_248 ( );
FILL FILL_30_DFFSR_248 ( );
FILL FILL_31_DFFSR_248 ( );
FILL FILL_32_DFFSR_248 ( );
FILL FILL_33_DFFSR_248 ( );
FILL FILL_34_DFFSR_248 ( );
FILL FILL_35_DFFSR_248 ( );
FILL FILL_36_DFFSR_248 ( );
FILL FILL_37_DFFSR_248 ( );
FILL FILL_38_DFFSR_248 ( );
FILL FILL_39_DFFSR_248 ( );
FILL FILL_40_DFFSR_248 ( );
FILL FILL_41_DFFSR_248 ( );
FILL FILL_42_DFFSR_248 ( );
FILL FILL_43_DFFSR_248 ( );
FILL FILL_44_DFFSR_248 ( );
FILL FILL_45_DFFSR_248 ( );
FILL FILL_46_DFFSR_248 ( );
FILL FILL_47_DFFSR_248 ( );
FILL FILL_48_DFFSR_248 ( );
FILL FILL_49_DFFSR_248 ( );
FILL FILL_50_DFFSR_248 ( );
FILL FILL_51_DFFSR_248 ( );
FILL FILL_0_INVX1_179 ( );
FILL FILL_1_INVX1_179 ( );
FILL FILL_2_INVX1_179 ( );
FILL FILL_3_INVX1_179 ( );
FILL FILL_4_INVX1_179 ( );
FILL FILL_0_NAND3X1_241 ( );
FILL FILL_1_NAND3X1_241 ( );
FILL FILL_2_NAND3X1_241 ( );
FILL FILL_3_NAND3X1_241 ( );
FILL FILL_4_NAND3X1_241 ( );
FILL FILL_5_NAND3X1_241 ( );
FILL FILL_6_NAND3X1_241 ( );
FILL FILL_7_NAND3X1_241 ( );
FILL FILL_8_NAND3X1_241 ( );
FILL FILL_9_NAND3X1_241 ( );
FILL FILL_0_AOI21X1_39 ( );
FILL FILL_1_AOI21X1_39 ( );
FILL FILL_2_AOI21X1_39 ( );
FILL FILL_3_AOI21X1_39 ( );
FILL FILL_4_AOI21X1_39 ( );
FILL FILL_5_AOI21X1_39 ( );
FILL FILL_6_AOI21X1_39 ( );
FILL FILL_7_AOI21X1_39 ( );
FILL FILL_8_AOI21X1_39 ( );
FILL FILL_0_NAND2X1_111 ( );
FILL FILL_1_NAND2X1_111 ( );
FILL FILL_2_NAND2X1_111 ( );
FILL FILL_3_NAND2X1_111 ( );
FILL FILL_4_NAND2X1_111 ( );
FILL FILL_5_NAND2X1_111 ( );
FILL FILL_6_NAND2X1_111 ( );
FILL FILL_0_OAI21X1_79 ( );
FILL FILL_1_OAI21X1_79 ( );
FILL FILL_2_OAI21X1_79 ( );
FILL FILL_3_OAI21X1_79 ( );
FILL FILL_4_OAI21X1_79 ( );
FILL FILL_5_OAI21X1_79 ( );
FILL FILL_6_OAI21X1_79 ( );
FILL FILL_7_OAI21X1_79 ( );
FILL FILL_8_OAI21X1_79 ( );
FILL FILL_0_OAI21X1_77 ( );
FILL FILL_1_OAI21X1_77 ( );
FILL FILL_2_OAI21X1_77 ( );
FILL FILL_3_OAI21X1_77 ( );
FILL FILL_4_OAI21X1_77 ( );
FILL FILL_5_OAI21X1_77 ( );
FILL FILL_6_OAI21X1_77 ( );
FILL FILL_7_OAI21X1_77 ( );
FILL FILL_8_OAI21X1_77 ( );
FILL FILL_0_DFFSR_8 ( );
FILL FILL_1_DFFSR_8 ( );
FILL FILL_2_DFFSR_8 ( );
FILL FILL_3_DFFSR_8 ( );
FILL FILL_4_DFFSR_8 ( );
FILL FILL_5_DFFSR_8 ( );
FILL FILL_6_DFFSR_8 ( );
FILL FILL_7_DFFSR_8 ( );
FILL FILL_8_DFFSR_8 ( );
FILL FILL_9_DFFSR_8 ( );
FILL FILL_10_DFFSR_8 ( );
FILL FILL_11_DFFSR_8 ( );
FILL FILL_12_DFFSR_8 ( );
FILL FILL_13_DFFSR_8 ( );
FILL FILL_14_DFFSR_8 ( );
FILL FILL_15_DFFSR_8 ( );
FILL FILL_16_DFFSR_8 ( );
FILL FILL_17_DFFSR_8 ( );
FILL FILL_18_DFFSR_8 ( );
FILL FILL_19_DFFSR_8 ( );
FILL FILL_20_DFFSR_8 ( );
FILL FILL_21_DFFSR_8 ( );
FILL FILL_22_DFFSR_8 ( );
FILL FILL_23_DFFSR_8 ( );
FILL FILL_24_DFFSR_8 ( );
FILL FILL_25_DFFSR_8 ( );
FILL FILL_26_DFFSR_8 ( );
FILL FILL_27_DFFSR_8 ( );
FILL FILL_28_DFFSR_8 ( );
FILL FILL_29_DFFSR_8 ( );
FILL FILL_30_DFFSR_8 ( );
FILL FILL_31_DFFSR_8 ( );
FILL FILL_32_DFFSR_8 ( );
FILL FILL_33_DFFSR_8 ( );
FILL FILL_34_DFFSR_8 ( );
FILL FILL_35_DFFSR_8 ( );
FILL FILL_36_DFFSR_8 ( );
FILL FILL_37_DFFSR_8 ( );
FILL FILL_38_DFFSR_8 ( );
FILL FILL_39_DFFSR_8 ( );
FILL FILL_40_DFFSR_8 ( );
FILL FILL_41_DFFSR_8 ( );
FILL FILL_42_DFFSR_8 ( );
FILL FILL_43_DFFSR_8 ( );
FILL FILL_44_DFFSR_8 ( );
FILL FILL_45_DFFSR_8 ( );
FILL FILL_46_DFFSR_8 ( );
FILL FILL_47_DFFSR_8 ( );
FILL FILL_48_DFFSR_8 ( );
FILL FILL_49_DFFSR_8 ( );
FILL FILL_50_DFFSR_8 ( );
FILL FILL_51_DFFSR_8 ( );
FILL FILL_0_DFFSR_12 ( );
FILL FILL_1_DFFSR_12 ( );
FILL FILL_2_DFFSR_12 ( );
FILL FILL_3_DFFSR_12 ( );
FILL FILL_4_DFFSR_12 ( );
FILL FILL_5_DFFSR_12 ( );
FILL FILL_6_DFFSR_12 ( );
FILL FILL_7_DFFSR_12 ( );
FILL FILL_8_DFFSR_12 ( );
FILL FILL_9_DFFSR_12 ( );
FILL FILL_10_DFFSR_12 ( );
FILL FILL_11_DFFSR_12 ( );
FILL FILL_12_DFFSR_12 ( );
FILL FILL_13_DFFSR_12 ( );
FILL FILL_14_DFFSR_12 ( );
FILL FILL_15_DFFSR_12 ( );
FILL FILL_16_DFFSR_12 ( );
FILL FILL_17_DFFSR_12 ( );
FILL FILL_18_DFFSR_12 ( );
FILL FILL_19_DFFSR_12 ( );
FILL FILL_20_DFFSR_12 ( );
FILL FILL_21_DFFSR_12 ( );
FILL FILL_22_DFFSR_12 ( );
FILL FILL_23_DFFSR_12 ( );
FILL FILL_24_DFFSR_12 ( );
FILL FILL_25_DFFSR_12 ( );
FILL FILL_26_DFFSR_12 ( );
FILL FILL_27_DFFSR_12 ( );
FILL FILL_28_DFFSR_12 ( );
FILL FILL_29_DFFSR_12 ( );
FILL FILL_30_DFFSR_12 ( );
FILL FILL_31_DFFSR_12 ( );
FILL FILL_32_DFFSR_12 ( );
FILL FILL_33_DFFSR_12 ( );
FILL FILL_34_DFFSR_12 ( );
FILL FILL_35_DFFSR_12 ( );
FILL FILL_36_DFFSR_12 ( );
FILL FILL_37_DFFSR_12 ( );
FILL FILL_38_DFFSR_12 ( );
FILL FILL_39_DFFSR_12 ( );
FILL FILL_40_DFFSR_12 ( );
FILL FILL_41_DFFSR_12 ( );
FILL FILL_42_DFFSR_12 ( );
FILL FILL_43_DFFSR_12 ( );
FILL FILL_44_DFFSR_12 ( );
FILL FILL_45_DFFSR_12 ( );
FILL FILL_46_DFFSR_12 ( );
FILL FILL_47_DFFSR_12 ( );
FILL FILL_48_DFFSR_12 ( );
FILL FILL_49_DFFSR_12 ( );
FILL FILL_50_DFFSR_12 ( );
FILL FILL_0_NAND3X1_25 ( );
FILL FILL_1_NAND3X1_25 ( );
FILL FILL_2_NAND3X1_25 ( );
FILL FILL_3_NAND3X1_25 ( );
FILL FILL_4_NAND3X1_25 ( );
FILL FILL_5_NAND3X1_25 ( );
FILL FILL_6_NAND3X1_25 ( );
FILL FILL_7_NAND3X1_25 ( );
FILL FILL_8_NAND3X1_25 ( );
FILL FILL_0_NAND3X1_28 ( );
FILL FILL_1_NAND3X1_28 ( );
FILL FILL_2_NAND3X1_28 ( );
FILL FILL_3_NAND3X1_28 ( );
FILL FILL_4_NAND3X1_28 ( );
FILL FILL_5_NAND3X1_28 ( );
FILL FILL_6_NAND3X1_28 ( );
FILL FILL_7_NAND3X1_28 ( );
FILL FILL_8_NAND3X1_28 ( );
FILL FILL_0_NAND2X1_26 ( );
FILL FILL_1_NAND2X1_26 ( );
FILL FILL_2_NAND2X1_26 ( );
FILL FILL_3_NAND2X1_26 ( );
FILL FILL_4_NAND2X1_26 ( );
FILL FILL_5_NAND2X1_26 ( );
FILL FILL_6_NAND2X1_26 ( );
FILL FILL_0_NAND3X1_60 ( );
FILL FILL_1_NAND3X1_60 ( );
FILL FILL_2_NAND3X1_60 ( );
FILL FILL_3_NAND3X1_60 ( );
FILL FILL_4_NAND3X1_60 ( );
FILL FILL_5_NAND3X1_60 ( );
FILL FILL_6_NAND3X1_60 ( );
FILL FILL_7_NAND3X1_60 ( );
FILL FILL_8_NAND3X1_60 ( );
FILL FILL_0_BUFX2_17 ( );
FILL FILL_1_BUFX2_17 ( );
FILL FILL_2_BUFX2_17 ( );
FILL FILL_3_BUFX2_17 ( );
FILL FILL_4_BUFX2_17 ( );
FILL FILL_5_BUFX2_17 ( );
FILL FILL_6_BUFX2_17 ( );
FILL FILL_0_AND2X2_5 ( );
FILL FILL_1_AND2X2_5 ( );
FILL FILL_2_AND2X2_5 ( );
FILL FILL_3_AND2X2_5 ( );
FILL FILL_4_AND2X2_5 ( );
FILL FILL_5_AND2X2_5 ( );
FILL FILL_6_AND2X2_5 ( );
FILL FILL_7_AND2X2_5 ( );
FILL FILL_8_AND2X2_5 ( );
FILL FILL_0_BUFX2_15 ( );
FILL FILL_1_BUFX2_15 ( );
FILL FILL_2_BUFX2_15 ( );
FILL FILL_3_BUFX2_15 ( );
FILL FILL_4_BUFX2_15 ( );
FILL FILL_5_BUFX2_15 ( );
FILL FILL_6_BUFX2_15 ( );
FILL FILL_0_INVX1_52 ( );
FILL FILL_1_INVX1_52 ( );
FILL FILL_2_INVX1_52 ( );
FILL FILL_3_INVX1_52 ( );
FILL FILL_4_INVX1_52 ( );
FILL FILL_0_OAI21X1_7 ( );
FILL FILL_1_OAI21X1_7 ( );
FILL FILL_2_OAI21X1_7 ( );
FILL FILL_3_OAI21X1_7 ( );
FILL FILL_4_OAI21X1_7 ( );
FILL FILL_5_OAI21X1_7 ( );
FILL FILL_6_OAI21X1_7 ( );
FILL FILL_7_OAI21X1_7 ( );
FILL FILL_8_OAI21X1_7 ( );
FILL FILL_9_OAI21X1_7 ( );
FILL FILL_0_NAND2X1_23 ( );
FILL FILL_1_NAND2X1_23 ( );
FILL FILL_2_NAND2X1_23 ( );
FILL FILL_3_NAND2X1_23 ( );
FILL FILL_4_NAND2X1_23 ( );
FILL FILL_5_NAND2X1_23 ( );
FILL FILL_6_NAND2X1_23 ( );
FILL FILL_0_AOI22X1_7 ( );
FILL FILL_1_AOI22X1_7 ( );
FILL FILL_2_AOI22X1_7 ( );
FILL FILL_3_AOI22X1_7 ( );
FILL FILL_4_AOI22X1_7 ( );
FILL FILL_5_AOI22X1_7 ( );
FILL FILL_6_AOI22X1_7 ( );
FILL FILL_7_AOI22X1_7 ( );
FILL FILL_8_AOI22X1_7 ( );
FILL FILL_9_AOI22X1_7 ( );
FILL FILL_10_AOI22X1_7 ( );
FILL FILL_11_AOI22X1_7 ( );
FILL FILL_0_DFFSR_111 ( );
FILL FILL_1_DFFSR_111 ( );
FILL FILL_2_DFFSR_111 ( );
FILL FILL_3_DFFSR_111 ( );
FILL FILL_4_DFFSR_111 ( );
FILL FILL_5_DFFSR_111 ( );
FILL FILL_6_DFFSR_111 ( );
FILL FILL_7_DFFSR_111 ( );
FILL FILL_8_DFFSR_111 ( );
FILL FILL_9_DFFSR_111 ( );
FILL FILL_10_DFFSR_111 ( );
FILL FILL_11_DFFSR_111 ( );
FILL FILL_12_DFFSR_111 ( );
FILL FILL_13_DFFSR_111 ( );
FILL FILL_14_DFFSR_111 ( );
FILL FILL_15_DFFSR_111 ( );
FILL FILL_16_DFFSR_111 ( );
FILL FILL_17_DFFSR_111 ( );
FILL FILL_18_DFFSR_111 ( );
FILL FILL_19_DFFSR_111 ( );
FILL FILL_20_DFFSR_111 ( );
FILL FILL_21_DFFSR_111 ( );
FILL FILL_22_DFFSR_111 ( );
FILL FILL_23_DFFSR_111 ( );
FILL FILL_24_DFFSR_111 ( );
FILL FILL_25_DFFSR_111 ( );
FILL FILL_26_DFFSR_111 ( );
FILL FILL_27_DFFSR_111 ( );
FILL FILL_28_DFFSR_111 ( );
FILL FILL_29_DFFSR_111 ( );
FILL FILL_30_DFFSR_111 ( );
FILL FILL_31_DFFSR_111 ( );
FILL FILL_32_DFFSR_111 ( );
FILL FILL_33_DFFSR_111 ( );
FILL FILL_34_DFFSR_111 ( );
FILL FILL_35_DFFSR_111 ( );
FILL FILL_36_DFFSR_111 ( );
FILL FILL_37_DFFSR_111 ( );
FILL FILL_38_DFFSR_111 ( );
FILL FILL_39_DFFSR_111 ( );
FILL FILL_40_DFFSR_111 ( );
FILL FILL_41_DFFSR_111 ( );
FILL FILL_42_DFFSR_111 ( );
FILL FILL_43_DFFSR_111 ( );
FILL FILL_44_DFFSR_111 ( );
FILL FILL_45_DFFSR_111 ( );
FILL FILL_46_DFFSR_111 ( );
FILL FILL_47_DFFSR_111 ( );
FILL FILL_48_DFFSR_111 ( );
FILL FILL_49_DFFSR_111 ( );
FILL FILL_50_DFFSR_111 ( );
FILL FILL_51_DFFSR_111 ( );
FILL FILL_0_NAND3X1_33 ( );
FILL FILL_1_NAND3X1_33 ( );
FILL FILL_2_NAND3X1_33 ( );
FILL FILL_3_NAND3X1_33 ( );
FILL FILL_4_NAND3X1_33 ( );
FILL FILL_5_NAND3X1_33 ( );
FILL FILL_6_NAND3X1_33 ( );
FILL FILL_7_NAND3X1_33 ( );
FILL FILL_8_NAND3X1_33 ( );
FILL FILL_9_NAND3X1_33 ( );
FILL FILL_0_NAND3X1_35 ( );
FILL FILL_1_NAND3X1_35 ( );
FILL FILL_2_NAND3X1_35 ( );
FILL FILL_3_NAND3X1_35 ( );
FILL FILL_4_NAND3X1_35 ( );
FILL FILL_5_NAND3X1_35 ( );
FILL FILL_6_NAND3X1_35 ( );
FILL FILL_7_NAND3X1_35 ( );
FILL FILL_8_NAND3X1_35 ( );
FILL FILL_0_AND2X2_10 ( );
FILL FILL_1_AND2X2_10 ( );
FILL FILL_2_AND2X2_10 ( );
FILL FILL_3_AND2X2_10 ( );
FILL FILL_4_AND2X2_10 ( );
FILL FILL_5_AND2X2_10 ( );
FILL FILL_6_AND2X2_10 ( );
FILL FILL_7_AND2X2_10 ( );
FILL FILL_8_AND2X2_10 ( );
FILL FILL_9_AND2X2_10 ( );
FILL FILL_0_NAND3X1_36 ( );
FILL FILL_1_NAND3X1_36 ( );
FILL FILL_2_NAND3X1_36 ( );
FILL FILL_3_NAND3X1_36 ( );
FILL FILL_4_NAND3X1_36 ( );
FILL FILL_5_NAND3X1_36 ( );
FILL FILL_6_NAND3X1_36 ( );
FILL FILL_7_NAND3X1_36 ( );
FILL FILL_8_NAND3X1_36 ( );
FILL FILL_0_NAND2X1_20 ( );
FILL FILL_1_NAND2X1_20 ( );
FILL FILL_2_NAND2X1_20 ( );
FILL FILL_3_NAND2X1_20 ( );
FILL FILL_4_NAND2X1_20 ( );
FILL FILL_5_NAND2X1_20 ( );
FILL FILL_6_NAND2X1_20 ( );
FILL FILL_0_OAI21X1_5 ( );
FILL FILL_1_OAI21X1_5 ( );
FILL FILL_2_OAI21X1_5 ( );
FILL FILL_3_OAI21X1_5 ( );
FILL FILL_4_OAI21X1_5 ( );
FILL FILL_5_OAI21X1_5 ( );
FILL FILL_6_OAI21X1_5 ( );
FILL FILL_7_OAI21X1_5 ( );
FILL FILL_8_OAI21X1_5 ( );
FILL FILL_0_NAND2X1_19 ( );
FILL FILL_1_NAND2X1_19 ( );
FILL FILL_2_NAND2X1_19 ( );
FILL FILL_3_NAND2X1_19 ( );
FILL FILL_4_NAND2X1_19 ( );
FILL FILL_5_NAND2X1_19 ( );
FILL FILL_6_NAND2X1_19 ( );
FILL FILL_0_DFFSR_85 ( );
FILL FILL_1_DFFSR_85 ( );
FILL FILL_2_DFFSR_85 ( );
FILL FILL_3_DFFSR_85 ( );
FILL FILL_4_DFFSR_85 ( );
FILL FILL_5_DFFSR_85 ( );
FILL FILL_6_DFFSR_85 ( );
FILL FILL_7_DFFSR_85 ( );
FILL FILL_8_DFFSR_85 ( );
FILL FILL_9_DFFSR_85 ( );
FILL FILL_10_DFFSR_85 ( );
FILL FILL_11_DFFSR_85 ( );
FILL FILL_12_DFFSR_85 ( );
FILL FILL_13_DFFSR_85 ( );
FILL FILL_14_DFFSR_85 ( );
FILL FILL_15_DFFSR_85 ( );
FILL FILL_16_DFFSR_85 ( );
FILL FILL_17_DFFSR_85 ( );
FILL FILL_18_DFFSR_85 ( );
FILL FILL_19_DFFSR_85 ( );
FILL FILL_20_DFFSR_85 ( );
FILL FILL_21_DFFSR_85 ( );
FILL FILL_22_DFFSR_85 ( );
FILL FILL_23_DFFSR_85 ( );
FILL FILL_24_DFFSR_85 ( );
FILL FILL_25_DFFSR_85 ( );
FILL FILL_26_DFFSR_85 ( );
FILL FILL_27_DFFSR_85 ( );
FILL FILL_28_DFFSR_85 ( );
FILL FILL_29_DFFSR_85 ( );
FILL FILL_30_DFFSR_85 ( );
FILL FILL_31_DFFSR_85 ( );
FILL FILL_32_DFFSR_85 ( );
FILL FILL_33_DFFSR_85 ( );
FILL FILL_34_DFFSR_85 ( );
FILL FILL_35_DFFSR_85 ( );
FILL FILL_36_DFFSR_85 ( );
FILL FILL_37_DFFSR_85 ( );
FILL FILL_38_DFFSR_85 ( );
FILL FILL_39_DFFSR_85 ( );
FILL FILL_40_DFFSR_85 ( );
FILL FILL_41_DFFSR_85 ( );
FILL FILL_42_DFFSR_85 ( );
FILL FILL_43_DFFSR_85 ( );
FILL FILL_44_DFFSR_85 ( );
FILL FILL_45_DFFSR_85 ( );
FILL FILL_46_DFFSR_85 ( );
FILL FILL_47_DFFSR_85 ( );
FILL FILL_48_DFFSR_85 ( );
FILL FILL_49_DFFSR_85 ( );
FILL FILL_50_DFFSR_85 ( );
FILL FILL_0_DFFSR_250 ( );
FILL FILL_1_DFFSR_250 ( );
FILL FILL_2_DFFSR_250 ( );
FILL FILL_3_DFFSR_250 ( );
FILL FILL_4_DFFSR_250 ( );
FILL FILL_5_DFFSR_250 ( );
FILL FILL_6_DFFSR_250 ( );
FILL FILL_7_DFFSR_250 ( );
FILL FILL_8_DFFSR_250 ( );
FILL FILL_9_DFFSR_250 ( );
FILL FILL_10_DFFSR_250 ( );
FILL FILL_11_DFFSR_250 ( );
FILL FILL_12_DFFSR_250 ( );
FILL FILL_13_DFFSR_250 ( );
FILL FILL_14_DFFSR_250 ( );
FILL FILL_15_DFFSR_250 ( );
FILL FILL_16_DFFSR_250 ( );
FILL FILL_17_DFFSR_250 ( );
FILL FILL_18_DFFSR_250 ( );
FILL FILL_19_DFFSR_250 ( );
FILL FILL_20_DFFSR_250 ( );
FILL FILL_21_DFFSR_250 ( );
FILL FILL_22_DFFSR_250 ( );
FILL FILL_23_DFFSR_250 ( );
FILL FILL_24_DFFSR_250 ( );
FILL FILL_25_DFFSR_250 ( );
FILL FILL_26_DFFSR_250 ( );
FILL FILL_27_DFFSR_250 ( );
FILL FILL_28_DFFSR_250 ( );
FILL FILL_29_DFFSR_250 ( );
FILL FILL_30_DFFSR_250 ( );
FILL FILL_31_DFFSR_250 ( );
FILL FILL_32_DFFSR_250 ( );
FILL FILL_33_DFFSR_250 ( );
FILL FILL_34_DFFSR_250 ( );
FILL FILL_35_DFFSR_250 ( );
FILL FILL_36_DFFSR_250 ( );
FILL FILL_37_DFFSR_250 ( );
FILL FILL_38_DFFSR_250 ( );
FILL FILL_39_DFFSR_250 ( );
FILL FILL_40_DFFSR_250 ( );
FILL FILL_41_DFFSR_250 ( );
FILL FILL_42_DFFSR_250 ( );
FILL FILL_43_DFFSR_250 ( );
FILL FILL_44_DFFSR_250 ( );
FILL FILL_45_DFFSR_250 ( );
FILL FILL_46_DFFSR_250 ( );
FILL FILL_47_DFFSR_250 ( );
FILL FILL_48_DFFSR_250 ( );
FILL FILL_49_DFFSR_250 ( );
FILL FILL_50_DFFSR_250 ( );
FILL FILL_0_CLKBUF1_1 ( );
FILL FILL_1_CLKBUF1_1 ( );
FILL FILL_2_CLKBUF1_1 ( );
FILL FILL_3_CLKBUF1_1 ( );
FILL FILL_4_CLKBUF1_1 ( );
FILL FILL_5_CLKBUF1_1 ( );
FILL FILL_6_CLKBUF1_1 ( );
FILL FILL_7_CLKBUF1_1 ( );
FILL FILL_8_CLKBUF1_1 ( );
FILL FILL_9_CLKBUF1_1 ( );
FILL FILL_10_CLKBUF1_1 ( );
FILL FILL_11_CLKBUF1_1 ( );
FILL FILL_12_CLKBUF1_1 ( );
FILL FILL_13_CLKBUF1_1 ( );
FILL FILL_14_CLKBUF1_1 ( );
FILL FILL_15_CLKBUF1_1 ( );
FILL FILL_16_CLKBUF1_1 ( );
FILL FILL_17_CLKBUF1_1 ( );
FILL FILL_18_CLKBUF1_1 ( );
FILL FILL_19_CLKBUF1_1 ( );
FILL FILL_20_CLKBUF1_1 ( );
FILL FILL_0_NAND3X1_239 ( );
FILL FILL_1_NAND3X1_239 ( );
FILL FILL_2_NAND3X1_239 ( );
FILL FILL_3_NAND3X1_239 ( );
FILL FILL_4_NAND3X1_239 ( );
FILL FILL_5_NAND3X1_239 ( );
FILL FILL_6_NAND3X1_239 ( );
FILL FILL_7_NAND3X1_239 ( );
FILL FILL_8_NAND3X1_239 ( );
FILL FILL_9_NAND3X1_239 ( );
FILL FILL_0_NAND3X1_240 ( );
FILL FILL_1_NAND3X1_240 ( );
FILL FILL_2_NAND3X1_240 ( );
FILL FILL_3_NAND3X1_240 ( );
FILL FILL_4_NAND3X1_240 ( );
FILL FILL_5_NAND3X1_240 ( );
FILL FILL_6_NAND3X1_240 ( );
FILL FILL_7_NAND3X1_240 ( );
FILL FILL_8_NAND3X1_240 ( );
FILL FILL_0_INVX1_176 ( );
FILL FILL_1_INVX1_176 ( );
FILL FILL_2_INVX1_176 ( );
FILL FILL_3_INVX1_176 ( );
FILL FILL_4_INVX1_176 ( );
FILL FILL_0_NAND2X1_108 ( );
FILL FILL_1_NAND2X1_108 ( );
FILL FILL_2_NAND2X1_108 ( );
FILL FILL_3_NAND2X1_108 ( );
FILL FILL_4_NAND2X1_108 ( );
FILL FILL_5_NAND2X1_108 ( );
FILL FILL_6_NAND2X1_108 ( );
FILL FILL_0_NOR2X1_72 ( );
FILL FILL_1_NOR2X1_72 ( );
FILL FILL_2_NOR2X1_72 ( );
FILL FILL_3_NOR2X1_72 ( );
FILL FILL_4_NOR2X1_72 ( );
FILL FILL_5_NOR2X1_72 ( );
FILL FILL_6_NOR2X1_72 ( );
FILL FILL_0_DFFPOSX1_41 ( );
FILL FILL_1_DFFPOSX1_41 ( );
FILL FILL_2_DFFPOSX1_41 ( );
FILL FILL_3_DFFPOSX1_41 ( );
FILL FILL_4_DFFPOSX1_41 ( );
FILL FILL_5_DFFPOSX1_41 ( );
FILL FILL_6_DFFPOSX1_41 ( );
FILL FILL_7_DFFPOSX1_41 ( );
FILL FILL_8_DFFPOSX1_41 ( );
FILL FILL_9_DFFPOSX1_41 ( );
FILL FILL_10_DFFPOSX1_41 ( );
FILL FILL_11_DFFPOSX1_41 ( );
FILL FILL_12_DFFPOSX1_41 ( );
FILL FILL_13_DFFPOSX1_41 ( );
FILL FILL_14_DFFPOSX1_41 ( );
FILL FILL_15_DFFPOSX1_41 ( );
FILL FILL_16_DFFPOSX1_41 ( );
FILL FILL_17_DFFPOSX1_41 ( );
FILL FILL_18_DFFPOSX1_41 ( );
FILL FILL_19_DFFPOSX1_41 ( );
FILL FILL_20_DFFPOSX1_41 ( );
FILL FILL_21_DFFPOSX1_41 ( );
FILL FILL_22_DFFPOSX1_41 ( );
FILL FILL_23_DFFPOSX1_41 ( );
FILL FILL_24_DFFPOSX1_41 ( );
FILL FILL_25_DFFPOSX1_41 ( );
FILL FILL_26_DFFPOSX1_41 ( );
FILL FILL_27_DFFPOSX1_41 ( );
FILL FILL_0_AOI21X1_53 ( );
FILL FILL_1_AOI21X1_53 ( );
FILL FILL_2_AOI21X1_53 ( );
FILL FILL_3_AOI21X1_53 ( );
FILL FILL_4_AOI21X1_53 ( );
FILL FILL_5_AOI21X1_53 ( );
FILL FILL_6_AOI21X1_53 ( );
FILL FILL_7_AOI21X1_53 ( );
FILL FILL_8_AOI21X1_53 ( );
FILL FILL_9_AOI21X1_53 ( );
FILL FILL_0_CLKBUF1_37 ( );
FILL FILL_1_CLKBUF1_37 ( );
FILL FILL_2_CLKBUF1_37 ( );
FILL FILL_3_CLKBUF1_37 ( );
FILL FILL_4_CLKBUF1_37 ( );
FILL FILL_5_CLKBUF1_37 ( );
FILL FILL_6_CLKBUF1_37 ( );
FILL FILL_7_CLKBUF1_37 ( );
FILL FILL_8_CLKBUF1_37 ( );
FILL FILL_9_CLKBUF1_37 ( );
FILL FILL_10_CLKBUF1_37 ( );
FILL FILL_11_CLKBUF1_37 ( );
FILL FILL_12_CLKBUF1_37 ( );
FILL FILL_13_CLKBUF1_37 ( );
FILL FILL_14_CLKBUF1_37 ( );
FILL FILL_15_CLKBUF1_37 ( );
FILL FILL_16_CLKBUF1_37 ( );
FILL FILL_17_CLKBUF1_37 ( );
FILL FILL_18_CLKBUF1_37 ( );
FILL FILL_19_CLKBUF1_37 ( );
FILL FILL_20_CLKBUF1_37 ( );
FILL FILL_0_INVX1_25 ( );
FILL FILL_1_INVX1_25 ( );
FILL FILL_2_INVX1_25 ( );
FILL FILL_3_INVX1_25 ( );
FILL FILL_4_INVX1_25 ( );
FILL FILL_0_DFFSR_48 ( );
FILL FILL_1_DFFSR_48 ( );
FILL FILL_2_DFFSR_48 ( );
FILL FILL_3_DFFSR_48 ( );
FILL FILL_4_DFFSR_48 ( );
FILL FILL_5_DFFSR_48 ( );
FILL FILL_6_DFFSR_48 ( );
FILL FILL_7_DFFSR_48 ( );
FILL FILL_8_DFFSR_48 ( );
FILL FILL_9_DFFSR_48 ( );
FILL FILL_10_DFFSR_48 ( );
FILL FILL_11_DFFSR_48 ( );
FILL FILL_12_DFFSR_48 ( );
FILL FILL_13_DFFSR_48 ( );
FILL FILL_14_DFFSR_48 ( );
FILL FILL_15_DFFSR_48 ( );
FILL FILL_16_DFFSR_48 ( );
FILL FILL_17_DFFSR_48 ( );
FILL FILL_18_DFFSR_48 ( );
FILL FILL_19_DFFSR_48 ( );
FILL FILL_20_DFFSR_48 ( );
FILL FILL_21_DFFSR_48 ( );
FILL FILL_22_DFFSR_48 ( );
FILL FILL_23_DFFSR_48 ( );
FILL FILL_24_DFFSR_48 ( );
FILL FILL_25_DFFSR_48 ( );
FILL FILL_26_DFFSR_48 ( );
FILL FILL_27_DFFSR_48 ( );
FILL FILL_28_DFFSR_48 ( );
FILL FILL_29_DFFSR_48 ( );
FILL FILL_30_DFFSR_48 ( );
FILL FILL_31_DFFSR_48 ( );
FILL FILL_32_DFFSR_48 ( );
FILL FILL_33_DFFSR_48 ( );
FILL FILL_34_DFFSR_48 ( );
FILL FILL_35_DFFSR_48 ( );
FILL FILL_36_DFFSR_48 ( );
FILL FILL_37_DFFSR_48 ( );
FILL FILL_38_DFFSR_48 ( );
FILL FILL_39_DFFSR_48 ( );
FILL FILL_40_DFFSR_48 ( );
FILL FILL_41_DFFSR_48 ( );
FILL FILL_42_DFFSR_48 ( );
FILL FILL_43_DFFSR_48 ( );
FILL FILL_44_DFFSR_48 ( );
FILL FILL_45_DFFSR_48 ( );
FILL FILL_46_DFFSR_48 ( );
FILL FILL_47_DFFSR_48 ( );
FILL FILL_48_DFFSR_48 ( );
FILL FILL_49_DFFSR_48 ( );
FILL FILL_50_DFFSR_48 ( );
FILL FILL_51_DFFSR_48 ( );
FILL FILL_0_INVX1_24 ( );
FILL FILL_1_INVX1_24 ( );
FILL FILL_2_INVX1_24 ( );
FILL FILL_3_INVX1_24 ( );
FILL FILL_0_OAI22X1_10 ( );
FILL FILL_1_OAI22X1_10 ( );
FILL FILL_2_OAI22X1_10 ( );
FILL FILL_3_OAI22X1_10 ( );
FILL FILL_4_OAI22X1_10 ( );
FILL FILL_5_OAI22X1_10 ( );
FILL FILL_6_OAI22X1_10 ( );
FILL FILL_7_OAI22X1_10 ( );
FILL FILL_8_OAI22X1_10 ( );
FILL FILL_9_OAI22X1_10 ( );
FILL FILL_10_OAI22X1_10 ( );
FILL FILL_11_OAI22X1_10 ( );
FILL FILL_0_NAND3X1_57 ( );
FILL FILL_1_NAND3X1_57 ( );
FILL FILL_2_NAND3X1_57 ( );
FILL FILL_3_NAND3X1_57 ( );
FILL FILL_4_NAND3X1_57 ( );
FILL FILL_5_NAND3X1_57 ( );
FILL FILL_6_NAND3X1_57 ( );
FILL FILL_7_NAND3X1_57 ( );
FILL FILL_8_NAND3X1_57 ( );
FILL FILL_9_NAND3X1_57 ( );
FILL FILL_0_INVX1_53 ( );
FILL FILL_1_INVX1_53 ( );
FILL FILL_2_INVX1_53 ( );
FILL FILL_3_INVX1_53 ( );
FILL FILL_4_INVX1_53 ( );
FILL FILL_0_NAND3X1_49 ( );
FILL FILL_1_NAND3X1_49 ( );
FILL FILL_2_NAND3X1_49 ( );
FILL FILL_3_NAND3X1_49 ( );
FILL FILL_4_NAND3X1_49 ( );
FILL FILL_5_NAND3X1_49 ( );
FILL FILL_6_NAND3X1_49 ( );
FILL FILL_7_NAND3X1_49 ( );
FILL FILL_8_NAND3X1_49 ( );
FILL FILL_0_NAND3X1_52 ( );
FILL FILL_1_NAND3X1_52 ( );
FILL FILL_2_NAND3X1_52 ( );
FILL FILL_3_NAND3X1_52 ( );
FILL FILL_4_NAND3X1_52 ( );
FILL FILL_5_NAND3X1_52 ( );
FILL FILL_6_NAND3X1_52 ( );
FILL FILL_7_NAND3X1_52 ( );
FILL FILL_8_NAND3X1_52 ( );
FILL FILL_0_NOR2X1_26 ( );
FILL FILL_1_NOR2X1_26 ( );
FILL FILL_2_NOR2X1_26 ( );
FILL FILL_3_NOR2X1_26 ( );
FILL FILL_4_NOR2X1_26 ( );
FILL FILL_5_NOR2X1_26 ( );
FILL FILL_6_NOR2X1_26 ( );
FILL FILL_0_OAI22X1_22 ( );
FILL FILL_1_OAI22X1_22 ( );
FILL FILL_2_OAI22X1_22 ( );
FILL FILL_3_OAI22X1_22 ( );
FILL FILL_4_OAI22X1_22 ( );
FILL FILL_5_OAI22X1_22 ( );
FILL FILL_6_OAI22X1_22 ( );
FILL FILL_7_OAI22X1_22 ( );
FILL FILL_8_OAI22X1_22 ( );
FILL FILL_9_OAI22X1_22 ( );
FILL FILL_10_OAI22X1_22 ( );
FILL FILL_0_NOR2X1_11 ( );
FILL FILL_1_NOR2X1_11 ( );
FILL FILL_2_NOR2X1_11 ( );
FILL FILL_3_NOR2X1_11 ( );
FILL FILL_4_NOR2X1_11 ( );
FILL FILL_5_NOR2X1_11 ( );
FILL FILL_6_NOR2X1_11 ( );
FILL FILL_0_DFFSR_103 ( );
FILL FILL_1_DFFSR_103 ( );
FILL FILL_2_DFFSR_103 ( );
FILL FILL_3_DFFSR_103 ( );
FILL FILL_4_DFFSR_103 ( );
FILL FILL_5_DFFSR_103 ( );
FILL FILL_6_DFFSR_103 ( );
FILL FILL_7_DFFSR_103 ( );
FILL FILL_8_DFFSR_103 ( );
FILL FILL_9_DFFSR_103 ( );
FILL FILL_10_DFFSR_103 ( );
FILL FILL_11_DFFSR_103 ( );
FILL FILL_12_DFFSR_103 ( );
FILL FILL_13_DFFSR_103 ( );
FILL FILL_14_DFFSR_103 ( );
FILL FILL_15_DFFSR_103 ( );
FILL FILL_16_DFFSR_103 ( );
FILL FILL_17_DFFSR_103 ( );
FILL FILL_18_DFFSR_103 ( );
FILL FILL_19_DFFSR_103 ( );
FILL FILL_20_DFFSR_103 ( );
FILL FILL_21_DFFSR_103 ( );
FILL FILL_22_DFFSR_103 ( );
FILL FILL_23_DFFSR_103 ( );
FILL FILL_24_DFFSR_103 ( );
FILL FILL_25_DFFSR_103 ( );
FILL FILL_26_DFFSR_103 ( );
FILL FILL_27_DFFSR_103 ( );
FILL FILL_28_DFFSR_103 ( );
FILL FILL_29_DFFSR_103 ( );
FILL FILL_30_DFFSR_103 ( );
FILL FILL_31_DFFSR_103 ( );
FILL FILL_32_DFFSR_103 ( );
FILL FILL_33_DFFSR_103 ( );
FILL FILL_34_DFFSR_103 ( );
FILL FILL_35_DFFSR_103 ( );
FILL FILL_36_DFFSR_103 ( );
FILL FILL_37_DFFSR_103 ( );
FILL FILL_38_DFFSR_103 ( );
FILL FILL_39_DFFSR_103 ( );
FILL FILL_40_DFFSR_103 ( );
FILL FILL_41_DFFSR_103 ( );
FILL FILL_42_DFFSR_103 ( );
FILL FILL_43_DFFSR_103 ( );
FILL FILL_44_DFFSR_103 ( );
FILL FILL_45_DFFSR_103 ( );
FILL FILL_46_DFFSR_103 ( );
FILL FILL_47_DFFSR_103 ( );
FILL FILL_48_DFFSR_103 ( );
FILL FILL_49_DFFSR_103 ( );
FILL FILL_50_DFFSR_103 ( );
FILL FILL_0_NOR2X1_27 ( );
FILL FILL_1_NOR2X1_27 ( );
FILL FILL_2_NOR2X1_27 ( );
FILL FILL_3_NOR2X1_27 ( );
FILL FILL_4_NOR2X1_27 ( );
FILL FILL_5_NOR2X1_27 ( );
FILL FILL_6_NOR2X1_27 ( );
FILL FILL_0_NAND3X1_62 ( );
FILL FILL_1_NAND3X1_62 ( );
FILL FILL_2_NAND3X1_62 ( );
FILL FILL_3_NAND3X1_62 ( );
FILL FILL_4_NAND3X1_62 ( );
FILL FILL_5_NAND3X1_62 ( );
FILL FILL_6_NAND3X1_62 ( );
FILL FILL_7_NAND3X1_62 ( );
FILL FILL_8_NAND3X1_62 ( );
FILL FILL_9_NAND3X1_62 ( );
FILL FILL_0_NAND3X1_34 ( );
FILL FILL_1_NAND3X1_34 ( );
FILL FILL_2_NAND3X1_34 ( );
FILL FILL_3_NAND3X1_34 ( );
FILL FILL_4_NAND3X1_34 ( );
FILL FILL_5_NAND3X1_34 ( );
FILL FILL_6_NAND3X1_34 ( );
FILL FILL_7_NAND3X1_34 ( );
FILL FILL_8_NAND3X1_34 ( );
FILL FILL_0_DFFSR_45 ( );
FILL FILL_1_DFFSR_45 ( );
FILL FILL_2_DFFSR_45 ( );
FILL FILL_3_DFFSR_45 ( );
FILL FILL_4_DFFSR_45 ( );
FILL FILL_5_DFFSR_45 ( );
FILL FILL_6_DFFSR_45 ( );
FILL FILL_7_DFFSR_45 ( );
FILL FILL_8_DFFSR_45 ( );
FILL FILL_9_DFFSR_45 ( );
FILL FILL_10_DFFSR_45 ( );
FILL FILL_11_DFFSR_45 ( );
FILL FILL_12_DFFSR_45 ( );
FILL FILL_13_DFFSR_45 ( );
FILL FILL_14_DFFSR_45 ( );
FILL FILL_15_DFFSR_45 ( );
FILL FILL_16_DFFSR_45 ( );
FILL FILL_17_DFFSR_45 ( );
FILL FILL_18_DFFSR_45 ( );
FILL FILL_19_DFFSR_45 ( );
FILL FILL_20_DFFSR_45 ( );
FILL FILL_21_DFFSR_45 ( );
FILL FILL_22_DFFSR_45 ( );
FILL FILL_23_DFFSR_45 ( );
FILL FILL_24_DFFSR_45 ( );
FILL FILL_25_DFFSR_45 ( );
FILL FILL_26_DFFSR_45 ( );
FILL FILL_27_DFFSR_45 ( );
FILL FILL_28_DFFSR_45 ( );
FILL FILL_29_DFFSR_45 ( );
FILL FILL_30_DFFSR_45 ( );
FILL FILL_31_DFFSR_45 ( );
FILL FILL_32_DFFSR_45 ( );
FILL FILL_33_DFFSR_45 ( );
FILL FILL_34_DFFSR_45 ( );
FILL FILL_35_DFFSR_45 ( );
FILL FILL_36_DFFSR_45 ( );
FILL FILL_37_DFFSR_45 ( );
FILL FILL_38_DFFSR_45 ( );
FILL FILL_39_DFFSR_45 ( );
FILL FILL_40_DFFSR_45 ( );
FILL FILL_41_DFFSR_45 ( );
FILL FILL_42_DFFSR_45 ( );
FILL FILL_43_DFFSR_45 ( );
FILL FILL_44_DFFSR_45 ( );
FILL FILL_45_DFFSR_45 ( );
FILL FILL_46_DFFSR_45 ( );
FILL FILL_47_DFFSR_45 ( );
FILL FILL_48_DFFSR_45 ( );
FILL FILL_49_DFFSR_45 ( );
FILL FILL_50_DFFSR_45 ( );
FILL FILL_51_DFFSR_45 ( );
FILL FILL_0_AOI22X1_5 ( );
FILL FILL_1_AOI22X1_5 ( );
FILL FILL_2_AOI22X1_5 ( );
FILL FILL_3_AOI22X1_5 ( );
FILL FILL_4_AOI22X1_5 ( );
FILL FILL_5_AOI22X1_5 ( );
FILL FILL_6_AOI22X1_5 ( );
FILL FILL_7_AOI22X1_5 ( );
FILL FILL_8_AOI22X1_5 ( );
FILL FILL_9_AOI22X1_5 ( );
FILL FILL_10_AOI22X1_5 ( );
FILL FILL_0_DFFSR_37 ( );
FILL FILL_1_DFFSR_37 ( );
FILL FILL_2_DFFSR_37 ( );
FILL FILL_3_DFFSR_37 ( );
FILL FILL_4_DFFSR_37 ( );
FILL FILL_5_DFFSR_37 ( );
FILL FILL_6_DFFSR_37 ( );
FILL FILL_7_DFFSR_37 ( );
FILL FILL_8_DFFSR_37 ( );
FILL FILL_9_DFFSR_37 ( );
FILL FILL_10_DFFSR_37 ( );
FILL FILL_11_DFFSR_37 ( );
FILL FILL_12_DFFSR_37 ( );
FILL FILL_13_DFFSR_37 ( );
FILL FILL_14_DFFSR_37 ( );
FILL FILL_15_DFFSR_37 ( );
FILL FILL_16_DFFSR_37 ( );
FILL FILL_17_DFFSR_37 ( );
FILL FILL_18_DFFSR_37 ( );
FILL FILL_19_DFFSR_37 ( );
FILL FILL_20_DFFSR_37 ( );
FILL FILL_21_DFFSR_37 ( );
FILL FILL_22_DFFSR_37 ( );
FILL FILL_23_DFFSR_37 ( );
FILL FILL_24_DFFSR_37 ( );
FILL FILL_25_DFFSR_37 ( );
FILL FILL_26_DFFSR_37 ( );
FILL FILL_27_DFFSR_37 ( );
FILL FILL_28_DFFSR_37 ( );
FILL FILL_29_DFFSR_37 ( );
FILL FILL_30_DFFSR_37 ( );
FILL FILL_31_DFFSR_37 ( );
FILL FILL_32_DFFSR_37 ( );
FILL FILL_33_DFFSR_37 ( );
FILL FILL_34_DFFSR_37 ( );
FILL FILL_35_DFFSR_37 ( );
FILL FILL_36_DFFSR_37 ( );
FILL FILL_37_DFFSR_37 ( );
FILL FILL_38_DFFSR_37 ( );
FILL FILL_39_DFFSR_37 ( );
FILL FILL_40_DFFSR_37 ( );
FILL FILL_41_DFFSR_37 ( );
FILL FILL_42_DFFSR_37 ( );
FILL FILL_43_DFFSR_37 ( );
FILL FILL_44_DFFSR_37 ( );
FILL FILL_45_DFFSR_37 ( );
FILL FILL_46_DFFSR_37 ( );
FILL FILL_47_DFFSR_37 ( );
FILL FILL_48_DFFSR_37 ( );
FILL FILL_49_DFFSR_37 ( );
FILL FILL_50_DFFSR_37 ( );
FILL FILL_0_DFFSR_256 ( );
FILL FILL_1_DFFSR_256 ( );
FILL FILL_2_DFFSR_256 ( );
FILL FILL_3_DFFSR_256 ( );
FILL FILL_4_DFFSR_256 ( );
FILL FILL_5_DFFSR_256 ( );
FILL FILL_6_DFFSR_256 ( );
FILL FILL_7_DFFSR_256 ( );
FILL FILL_8_DFFSR_256 ( );
FILL FILL_9_DFFSR_256 ( );
FILL FILL_10_DFFSR_256 ( );
FILL FILL_11_DFFSR_256 ( );
FILL FILL_12_DFFSR_256 ( );
FILL FILL_13_DFFSR_256 ( );
FILL FILL_14_DFFSR_256 ( );
FILL FILL_15_DFFSR_256 ( );
FILL FILL_16_DFFSR_256 ( );
FILL FILL_17_DFFSR_256 ( );
FILL FILL_18_DFFSR_256 ( );
FILL FILL_19_DFFSR_256 ( );
FILL FILL_20_DFFSR_256 ( );
FILL FILL_21_DFFSR_256 ( );
FILL FILL_22_DFFSR_256 ( );
FILL FILL_23_DFFSR_256 ( );
FILL FILL_24_DFFSR_256 ( );
FILL FILL_25_DFFSR_256 ( );
FILL FILL_26_DFFSR_256 ( );
FILL FILL_27_DFFSR_256 ( );
FILL FILL_28_DFFSR_256 ( );
FILL FILL_29_DFFSR_256 ( );
FILL FILL_30_DFFSR_256 ( );
FILL FILL_31_DFFSR_256 ( );
FILL FILL_32_DFFSR_256 ( );
FILL FILL_33_DFFSR_256 ( );
FILL FILL_34_DFFSR_256 ( );
FILL FILL_35_DFFSR_256 ( );
FILL FILL_36_DFFSR_256 ( );
FILL FILL_37_DFFSR_256 ( );
FILL FILL_38_DFFSR_256 ( );
FILL FILL_39_DFFSR_256 ( );
FILL FILL_40_DFFSR_256 ( );
FILL FILL_41_DFFSR_256 ( );
FILL FILL_42_DFFSR_256 ( );
FILL FILL_43_DFFSR_256 ( );
FILL FILL_44_DFFSR_256 ( );
FILL FILL_45_DFFSR_256 ( );
FILL FILL_46_DFFSR_256 ( );
FILL FILL_47_DFFSR_256 ( );
FILL FILL_48_DFFSR_256 ( );
FILL FILL_49_DFFSR_256 ( );
FILL FILL_50_DFFSR_256 ( );
FILL FILL_0_BUFX2_65 ( );
FILL FILL_1_BUFX2_65 ( );
FILL FILL_2_BUFX2_65 ( );
FILL FILL_3_BUFX2_65 ( );
FILL FILL_4_BUFX2_65 ( );
FILL FILL_5_BUFX2_65 ( );
FILL FILL_6_BUFX2_65 ( );
FILL FILL_0_OAI21X1_80 ( );
FILL FILL_1_OAI21X1_80 ( );
FILL FILL_2_OAI21X1_80 ( );
FILL FILL_3_OAI21X1_80 ( );
FILL FILL_4_OAI21X1_80 ( );
FILL FILL_5_OAI21X1_80 ( );
FILL FILL_6_OAI21X1_80 ( );
FILL FILL_7_OAI21X1_80 ( );
FILL FILL_8_OAI21X1_80 ( );
FILL FILL_0_NAND3X1_237 ( );
FILL FILL_1_NAND3X1_237 ( );
FILL FILL_2_NAND3X1_237 ( );
FILL FILL_3_NAND3X1_237 ( );
FILL FILL_4_NAND3X1_237 ( );
FILL FILL_5_NAND3X1_237 ( );
FILL FILL_6_NAND3X1_237 ( );
FILL FILL_7_NAND3X1_237 ( );
FILL FILL_8_NAND3X1_237 ( );
FILL FILL_0_NOR2X1_73 ( );
FILL FILL_1_NOR2X1_73 ( );
FILL FILL_2_NOR2X1_73 ( );
FILL FILL_3_NOR2X1_73 ( );
FILL FILL_4_NOR2X1_73 ( );
FILL FILL_5_NOR2X1_73 ( );
FILL FILL_6_NOR2X1_73 ( );
FILL FILL_0_NAND3X1_226 ( );
FILL FILL_1_NAND3X1_226 ( );
FILL FILL_2_NAND3X1_226 ( );
FILL FILL_3_NAND3X1_226 ( );
FILL FILL_4_NAND3X1_226 ( );
FILL FILL_5_NAND3X1_226 ( );
FILL FILL_6_NAND3X1_226 ( );
FILL FILL_7_NAND3X1_226 ( );
FILL FILL_8_NAND3X1_226 ( );
FILL FILL_0_NAND2X1_107 ( );
FILL FILL_1_NAND2X1_107 ( );
FILL FILL_2_NAND2X1_107 ( );
FILL FILL_3_NAND2X1_107 ( );
FILL FILL_4_NAND2X1_107 ( );
FILL FILL_5_NAND2X1_107 ( );
FILL FILL_6_NAND2X1_107 ( );
FILL FILL_0_INVX1_177 ( );
FILL FILL_1_INVX1_177 ( );
FILL FILL_2_INVX1_177 ( );
FILL FILL_3_INVX1_177 ( );
FILL FILL_0_CLKBUF1_4 ( );
FILL FILL_1_CLKBUF1_4 ( );
FILL FILL_2_CLKBUF1_4 ( );
FILL FILL_3_CLKBUF1_4 ( );
FILL FILL_4_CLKBUF1_4 ( );
FILL FILL_5_CLKBUF1_4 ( );
FILL FILL_6_CLKBUF1_4 ( );
FILL FILL_7_CLKBUF1_4 ( );
FILL FILL_8_CLKBUF1_4 ( );
FILL FILL_9_CLKBUF1_4 ( );
FILL FILL_10_CLKBUF1_4 ( );
FILL FILL_11_CLKBUF1_4 ( );
FILL FILL_12_CLKBUF1_4 ( );
FILL FILL_13_CLKBUF1_4 ( );
FILL FILL_14_CLKBUF1_4 ( );
FILL FILL_15_CLKBUF1_4 ( );
FILL FILL_16_CLKBUF1_4 ( );
FILL FILL_17_CLKBUF1_4 ( );
FILL FILL_18_CLKBUF1_4 ( );
FILL FILL_19_CLKBUF1_4 ( );
FILL FILL_0_DFFSR_60 ( );
FILL FILL_1_DFFSR_60 ( );
FILL FILL_2_DFFSR_60 ( );
FILL FILL_3_DFFSR_60 ( );
FILL FILL_4_DFFSR_60 ( );
FILL FILL_5_DFFSR_60 ( );
FILL FILL_6_DFFSR_60 ( );
FILL FILL_7_DFFSR_60 ( );
FILL FILL_8_DFFSR_60 ( );
FILL FILL_9_DFFSR_60 ( );
FILL FILL_10_DFFSR_60 ( );
FILL FILL_11_DFFSR_60 ( );
FILL FILL_12_DFFSR_60 ( );
FILL FILL_13_DFFSR_60 ( );
FILL FILL_14_DFFSR_60 ( );
FILL FILL_15_DFFSR_60 ( );
FILL FILL_16_DFFSR_60 ( );
FILL FILL_17_DFFSR_60 ( );
FILL FILL_18_DFFSR_60 ( );
FILL FILL_19_DFFSR_60 ( );
FILL FILL_20_DFFSR_60 ( );
FILL FILL_21_DFFSR_60 ( );
FILL FILL_22_DFFSR_60 ( );
FILL FILL_23_DFFSR_60 ( );
FILL FILL_24_DFFSR_60 ( );
FILL FILL_25_DFFSR_60 ( );
FILL FILL_26_DFFSR_60 ( );
FILL FILL_27_DFFSR_60 ( );
FILL FILL_28_DFFSR_60 ( );
FILL FILL_29_DFFSR_60 ( );
FILL FILL_30_DFFSR_60 ( );
FILL FILL_31_DFFSR_60 ( );
FILL FILL_32_DFFSR_60 ( );
FILL FILL_33_DFFSR_60 ( );
FILL FILL_34_DFFSR_60 ( );
FILL FILL_35_DFFSR_60 ( );
FILL FILL_36_DFFSR_60 ( );
FILL FILL_37_DFFSR_60 ( );
FILL FILL_38_DFFSR_60 ( );
FILL FILL_39_DFFSR_60 ( );
FILL FILL_40_DFFSR_60 ( );
FILL FILL_41_DFFSR_60 ( );
FILL FILL_42_DFFSR_60 ( );
FILL FILL_43_DFFSR_60 ( );
FILL FILL_44_DFFSR_60 ( );
FILL FILL_45_DFFSR_60 ( );
FILL FILL_46_DFFSR_60 ( );
FILL FILL_47_DFFSR_60 ( );
FILL FILL_48_DFFSR_60 ( );
FILL FILL_49_DFFSR_60 ( );
FILL FILL_50_DFFSR_60 ( );
FILL FILL_51_DFFSR_60 ( );
FILL FILL_0_DFFSR_64 ( );
FILL FILL_1_DFFSR_64 ( );
FILL FILL_2_DFFSR_64 ( );
FILL FILL_3_DFFSR_64 ( );
FILL FILL_4_DFFSR_64 ( );
FILL FILL_5_DFFSR_64 ( );
FILL FILL_6_DFFSR_64 ( );
FILL FILL_7_DFFSR_64 ( );
FILL FILL_8_DFFSR_64 ( );
FILL FILL_9_DFFSR_64 ( );
FILL FILL_10_DFFSR_64 ( );
FILL FILL_11_DFFSR_64 ( );
FILL FILL_12_DFFSR_64 ( );
FILL FILL_13_DFFSR_64 ( );
FILL FILL_14_DFFSR_64 ( );
FILL FILL_15_DFFSR_64 ( );
FILL FILL_16_DFFSR_64 ( );
FILL FILL_17_DFFSR_64 ( );
FILL FILL_18_DFFSR_64 ( );
FILL FILL_19_DFFSR_64 ( );
FILL FILL_20_DFFSR_64 ( );
FILL FILL_21_DFFSR_64 ( );
FILL FILL_22_DFFSR_64 ( );
FILL FILL_23_DFFSR_64 ( );
FILL FILL_24_DFFSR_64 ( );
FILL FILL_25_DFFSR_64 ( );
FILL FILL_26_DFFSR_64 ( );
FILL FILL_27_DFFSR_64 ( );
FILL FILL_28_DFFSR_64 ( );
FILL FILL_29_DFFSR_64 ( );
FILL FILL_30_DFFSR_64 ( );
FILL FILL_31_DFFSR_64 ( );
FILL FILL_32_DFFSR_64 ( );
FILL FILL_33_DFFSR_64 ( );
FILL FILL_34_DFFSR_64 ( );
FILL FILL_35_DFFSR_64 ( );
FILL FILL_36_DFFSR_64 ( );
FILL FILL_37_DFFSR_64 ( );
FILL FILL_38_DFFSR_64 ( );
FILL FILL_39_DFFSR_64 ( );
FILL FILL_40_DFFSR_64 ( );
FILL FILL_41_DFFSR_64 ( );
FILL FILL_42_DFFSR_64 ( );
FILL FILL_43_DFFSR_64 ( );
FILL FILL_44_DFFSR_64 ( );
FILL FILL_45_DFFSR_64 ( );
FILL FILL_46_DFFSR_64 ( );
FILL FILL_47_DFFSR_64 ( );
FILL FILL_48_DFFSR_64 ( );
FILL FILL_49_DFFSR_64 ( );
FILL FILL_50_DFFSR_64 ( );
FILL FILL_0_NAND2X1_18 ( );
FILL FILL_1_NAND2X1_18 ( );
FILL FILL_2_NAND2X1_18 ( );
FILL FILL_3_NAND2X1_18 ( );
FILL FILL_4_NAND2X1_18 ( );
FILL FILL_5_NAND2X1_18 ( );
FILL FILL_6_NAND2X1_18 ( );
FILL FILL_0_OAI22X1_19 ( );
FILL FILL_1_OAI22X1_19 ( );
FILL FILL_2_OAI22X1_19 ( );
FILL FILL_3_OAI22X1_19 ( );
FILL FILL_4_OAI22X1_19 ( );
FILL FILL_5_OAI22X1_19 ( );
FILL FILL_6_OAI22X1_19 ( );
FILL FILL_7_OAI22X1_19 ( );
FILL FILL_8_OAI22X1_19 ( );
FILL FILL_9_OAI22X1_19 ( );
FILL FILL_10_OAI22X1_19 ( );
FILL FILL_11_OAI22X1_19 ( );
FILL FILL_0_BUFX2_47 ( );
FILL FILL_1_BUFX2_47 ( );
FILL FILL_2_BUFX2_47 ( );
FILL FILL_3_BUFX2_47 ( );
FILL FILL_4_BUFX2_47 ( );
FILL FILL_5_BUFX2_47 ( );
FILL FILL_6_BUFX2_47 ( );
FILL FILL_0_NAND3X1_53 ( );
FILL FILL_1_NAND3X1_53 ( );
FILL FILL_2_NAND3X1_53 ( );
FILL FILL_3_NAND3X1_53 ( );
FILL FILL_4_NAND3X1_53 ( );
FILL FILL_5_NAND3X1_53 ( );
FILL FILL_6_NAND3X1_53 ( );
FILL FILL_7_NAND3X1_53 ( );
FILL FILL_8_NAND3X1_53 ( );
FILL FILL_9_NAND3X1_53 ( );
FILL FILL_0_NAND3X1_55 ( );
FILL FILL_1_NAND3X1_55 ( );
FILL FILL_2_NAND3X1_55 ( );
FILL FILL_3_NAND3X1_55 ( );
FILL FILL_4_NAND3X1_55 ( );
FILL FILL_5_NAND3X1_55 ( );
FILL FILL_6_NAND3X1_55 ( );
FILL FILL_7_NAND3X1_55 ( );
FILL FILL_8_NAND3X1_55 ( );
FILL FILL_0_NAND3X1_54 ( );
FILL FILL_1_NAND3X1_54 ( );
FILL FILL_2_NAND3X1_54 ( );
FILL FILL_3_NAND3X1_54 ( );
FILL FILL_4_NAND3X1_54 ( );
FILL FILL_5_NAND3X1_54 ( );
FILL FILL_6_NAND3X1_54 ( );
FILL FILL_7_NAND3X1_54 ( );
FILL FILL_8_NAND3X1_54 ( );
FILL FILL_0_CLKBUF1_38 ( );
FILL FILL_1_CLKBUF1_38 ( );
FILL FILL_2_CLKBUF1_38 ( );
FILL FILL_3_CLKBUF1_38 ( );
FILL FILL_4_CLKBUF1_38 ( );
FILL FILL_5_CLKBUF1_38 ( );
FILL FILL_6_CLKBUF1_38 ( );
FILL FILL_7_CLKBUF1_38 ( );
FILL FILL_8_CLKBUF1_38 ( );
FILL FILL_9_CLKBUF1_38 ( );
FILL FILL_10_CLKBUF1_38 ( );
FILL FILL_11_CLKBUF1_38 ( );
FILL FILL_12_CLKBUF1_38 ( );
FILL FILL_13_CLKBUF1_38 ( );
FILL FILL_14_CLKBUF1_38 ( );
FILL FILL_15_CLKBUF1_38 ( );
FILL FILL_16_CLKBUF1_38 ( );
FILL FILL_17_CLKBUF1_38 ( );
FILL FILL_18_CLKBUF1_38 ( );
FILL FILL_19_CLKBUF1_38 ( );
FILL FILL_20_CLKBUF1_38 ( );
FILL FILL_0_NAND3X1_45 ( );
FILL FILL_1_NAND3X1_45 ( );
FILL FILL_2_NAND3X1_45 ( );
FILL FILL_3_NAND3X1_45 ( );
FILL FILL_4_NAND3X1_45 ( );
FILL FILL_5_NAND3X1_45 ( );
FILL FILL_6_NAND3X1_45 ( );
FILL FILL_7_NAND3X1_45 ( );
FILL FILL_8_NAND3X1_45 ( );
FILL FILL_0_DFFSR_72 ( );
FILL FILL_1_DFFSR_72 ( );
FILL FILL_2_DFFSR_72 ( );
FILL FILL_3_DFFSR_72 ( );
FILL FILL_4_DFFSR_72 ( );
FILL FILL_5_DFFSR_72 ( );
FILL FILL_6_DFFSR_72 ( );
FILL FILL_7_DFFSR_72 ( );
FILL FILL_8_DFFSR_72 ( );
FILL FILL_9_DFFSR_72 ( );
FILL FILL_10_DFFSR_72 ( );
FILL FILL_11_DFFSR_72 ( );
FILL FILL_12_DFFSR_72 ( );
FILL FILL_13_DFFSR_72 ( );
FILL FILL_14_DFFSR_72 ( );
FILL FILL_15_DFFSR_72 ( );
FILL FILL_16_DFFSR_72 ( );
FILL FILL_17_DFFSR_72 ( );
FILL FILL_18_DFFSR_72 ( );
FILL FILL_19_DFFSR_72 ( );
FILL FILL_20_DFFSR_72 ( );
FILL FILL_21_DFFSR_72 ( );
FILL FILL_22_DFFSR_72 ( );
FILL FILL_23_DFFSR_72 ( );
FILL FILL_24_DFFSR_72 ( );
FILL FILL_25_DFFSR_72 ( );
FILL FILL_26_DFFSR_72 ( );
FILL FILL_27_DFFSR_72 ( );
FILL FILL_28_DFFSR_72 ( );
FILL FILL_29_DFFSR_72 ( );
FILL FILL_30_DFFSR_72 ( );
FILL FILL_31_DFFSR_72 ( );
FILL FILL_32_DFFSR_72 ( );
FILL FILL_33_DFFSR_72 ( );
FILL FILL_34_DFFSR_72 ( );
FILL FILL_35_DFFSR_72 ( );
FILL FILL_36_DFFSR_72 ( );
FILL FILL_37_DFFSR_72 ( );
FILL FILL_38_DFFSR_72 ( );
FILL FILL_39_DFFSR_72 ( );
FILL FILL_40_DFFSR_72 ( );
FILL FILL_41_DFFSR_72 ( );
FILL FILL_42_DFFSR_72 ( );
FILL FILL_43_DFFSR_72 ( );
FILL FILL_44_DFFSR_72 ( );
FILL FILL_45_DFFSR_72 ( );
FILL FILL_46_DFFSR_72 ( );
FILL FILL_47_DFFSR_72 ( );
FILL FILL_48_DFFSR_72 ( );
FILL FILL_49_DFFSR_72 ( );
FILL FILL_50_DFFSR_72 ( );
FILL FILL_51_DFFSR_72 ( );
FILL FILL_0_DFFSR_118 ( );
FILL FILL_1_DFFSR_118 ( );
FILL FILL_2_DFFSR_118 ( );
FILL FILL_3_DFFSR_118 ( );
FILL FILL_4_DFFSR_118 ( );
FILL FILL_5_DFFSR_118 ( );
FILL FILL_6_DFFSR_118 ( );
FILL FILL_7_DFFSR_118 ( );
FILL FILL_8_DFFSR_118 ( );
FILL FILL_9_DFFSR_118 ( );
FILL FILL_10_DFFSR_118 ( );
FILL FILL_11_DFFSR_118 ( );
FILL FILL_12_DFFSR_118 ( );
FILL FILL_13_DFFSR_118 ( );
FILL FILL_14_DFFSR_118 ( );
FILL FILL_15_DFFSR_118 ( );
FILL FILL_16_DFFSR_118 ( );
FILL FILL_17_DFFSR_118 ( );
FILL FILL_18_DFFSR_118 ( );
FILL FILL_19_DFFSR_118 ( );
FILL FILL_20_DFFSR_118 ( );
FILL FILL_21_DFFSR_118 ( );
FILL FILL_22_DFFSR_118 ( );
FILL FILL_23_DFFSR_118 ( );
FILL FILL_24_DFFSR_118 ( );
FILL FILL_25_DFFSR_118 ( );
FILL FILL_26_DFFSR_118 ( );
FILL FILL_27_DFFSR_118 ( );
FILL FILL_28_DFFSR_118 ( );
FILL FILL_29_DFFSR_118 ( );
FILL FILL_30_DFFSR_118 ( );
FILL FILL_31_DFFSR_118 ( );
FILL FILL_32_DFFSR_118 ( );
FILL FILL_33_DFFSR_118 ( );
FILL FILL_34_DFFSR_118 ( );
FILL FILL_35_DFFSR_118 ( );
FILL FILL_36_DFFSR_118 ( );
FILL FILL_37_DFFSR_118 ( );
FILL FILL_38_DFFSR_118 ( );
FILL FILL_39_DFFSR_118 ( );
FILL FILL_40_DFFSR_118 ( );
FILL FILL_41_DFFSR_118 ( );
FILL FILL_42_DFFSR_118 ( );
FILL FILL_43_DFFSR_118 ( );
FILL FILL_44_DFFSR_118 ( );
FILL FILL_45_DFFSR_118 ( );
FILL FILL_46_DFFSR_118 ( );
FILL FILL_47_DFFSR_118 ( );
FILL FILL_48_DFFSR_118 ( );
FILL FILL_49_DFFSR_118 ( );
FILL FILL_50_DFFSR_118 ( );
FILL FILL_0_DFFSR_93 ( );
FILL FILL_1_DFFSR_93 ( );
FILL FILL_2_DFFSR_93 ( );
FILL FILL_3_DFFSR_93 ( );
FILL FILL_4_DFFSR_93 ( );
FILL FILL_5_DFFSR_93 ( );
FILL FILL_6_DFFSR_93 ( );
FILL FILL_7_DFFSR_93 ( );
FILL FILL_8_DFFSR_93 ( );
FILL FILL_9_DFFSR_93 ( );
FILL FILL_10_DFFSR_93 ( );
FILL FILL_11_DFFSR_93 ( );
FILL FILL_12_DFFSR_93 ( );
FILL FILL_13_DFFSR_93 ( );
FILL FILL_14_DFFSR_93 ( );
FILL FILL_15_DFFSR_93 ( );
FILL FILL_16_DFFSR_93 ( );
FILL FILL_17_DFFSR_93 ( );
FILL FILL_18_DFFSR_93 ( );
FILL FILL_19_DFFSR_93 ( );
FILL FILL_20_DFFSR_93 ( );
FILL FILL_21_DFFSR_93 ( );
FILL FILL_22_DFFSR_93 ( );
FILL FILL_23_DFFSR_93 ( );
FILL FILL_24_DFFSR_93 ( );
FILL FILL_25_DFFSR_93 ( );
FILL FILL_26_DFFSR_93 ( );
FILL FILL_27_DFFSR_93 ( );
FILL FILL_28_DFFSR_93 ( );
FILL FILL_29_DFFSR_93 ( );
FILL FILL_30_DFFSR_93 ( );
FILL FILL_31_DFFSR_93 ( );
FILL FILL_32_DFFSR_93 ( );
FILL FILL_33_DFFSR_93 ( );
FILL FILL_34_DFFSR_93 ( );
FILL FILL_35_DFFSR_93 ( );
FILL FILL_36_DFFSR_93 ( );
FILL FILL_37_DFFSR_93 ( );
FILL FILL_38_DFFSR_93 ( );
FILL FILL_39_DFFSR_93 ( );
FILL FILL_40_DFFSR_93 ( );
FILL FILL_41_DFFSR_93 ( );
FILL FILL_42_DFFSR_93 ( );
FILL FILL_43_DFFSR_93 ( );
FILL FILL_44_DFFSR_93 ( );
FILL FILL_45_DFFSR_93 ( );
FILL FILL_46_DFFSR_93 ( );
FILL FILL_47_DFFSR_93 ( );
FILL FILL_48_DFFSR_93 ( );
FILL FILL_49_DFFSR_93 ( );
FILL FILL_50_DFFSR_93 ( );
FILL FILL_0_BUFX2_97 ( );
FILL FILL_1_BUFX2_97 ( );
FILL FILL_2_BUFX2_97 ( );
FILL FILL_3_BUFX2_97 ( );
FILL FILL_4_BUFX2_97 ( );
FILL FILL_5_BUFX2_97 ( );
FILL FILL_6_BUFX2_97 ( );
FILL FILL_0_DFFSR_242 ( );
FILL FILL_1_DFFSR_242 ( );
FILL FILL_2_DFFSR_242 ( );
FILL FILL_3_DFFSR_242 ( );
FILL FILL_4_DFFSR_242 ( );
FILL FILL_5_DFFSR_242 ( );
FILL FILL_6_DFFSR_242 ( );
FILL FILL_7_DFFSR_242 ( );
FILL FILL_8_DFFSR_242 ( );
FILL FILL_9_DFFSR_242 ( );
FILL FILL_10_DFFSR_242 ( );
FILL FILL_11_DFFSR_242 ( );
FILL FILL_12_DFFSR_242 ( );
FILL FILL_13_DFFSR_242 ( );
FILL FILL_14_DFFSR_242 ( );
FILL FILL_15_DFFSR_242 ( );
FILL FILL_16_DFFSR_242 ( );
FILL FILL_17_DFFSR_242 ( );
FILL FILL_18_DFFSR_242 ( );
FILL FILL_19_DFFSR_242 ( );
FILL FILL_20_DFFSR_242 ( );
FILL FILL_21_DFFSR_242 ( );
FILL FILL_22_DFFSR_242 ( );
FILL FILL_23_DFFSR_242 ( );
FILL FILL_24_DFFSR_242 ( );
FILL FILL_25_DFFSR_242 ( );
FILL FILL_26_DFFSR_242 ( );
FILL FILL_27_DFFSR_242 ( );
FILL FILL_28_DFFSR_242 ( );
FILL FILL_29_DFFSR_242 ( );
FILL FILL_30_DFFSR_242 ( );
FILL FILL_31_DFFSR_242 ( );
FILL FILL_32_DFFSR_242 ( );
FILL FILL_33_DFFSR_242 ( );
FILL FILL_34_DFFSR_242 ( );
FILL FILL_35_DFFSR_242 ( );
FILL FILL_36_DFFSR_242 ( );
FILL FILL_37_DFFSR_242 ( );
FILL FILL_38_DFFSR_242 ( );
FILL FILL_39_DFFSR_242 ( );
FILL FILL_40_DFFSR_242 ( );
FILL FILL_41_DFFSR_242 ( );
FILL FILL_42_DFFSR_242 ( );
FILL FILL_43_DFFSR_242 ( );
FILL FILL_44_DFFSR_242 ( );
FILL FILL_45_DFFSR_242 ( );
FILL FILL_46_DFFSR_242 ( );
FILL FILL_47_DFFSR_242 ( );
FILL FILL_48_DFFSR_242 ( );
FILL FILL_49_DFFSR_242 ( );
FILL FILL_50_DFFSR_242 ( );
FILL FILL_51_DFFSR_242 ( );
FILL FILL_0_OAI21X1_89 ( );
FILL FILL_1_OAI21X1_89 ( );
FILL FILL_2_OAI21X1_89 ( );
FILL FILL_3_OAI21X1_89 ( );
FILL FILL_4_OAI21X1_89 ( );
FILL FILL_5_OAI21X1_89 ( );
FILL FILL_6_OAI21X1_89 ( );
FILL FILL_7_OAI21X1_89 ( );
FILL FILL_8_OAI21X1_89 ( );
FILL FILL_0_OAI21X1_81 ( );
FILL FILL_1_OAI21X1_81 ( );
FILL FILL_2_OAI21X1_81 ( );
FILL FILL_3_OAI21X1_81 ( );
FILL FILL_4_OAI21X1_81 ( );
FILL FILL_5_OAI21X1_81 ( );
FILL FILL_6_OAI21X1_81 ( );
FILL FILL_7_OAI21X1_81 ( );
FILL FILL_8_OAI21X1_81 ( );
FILL FILL_9_OAI21X1_81 ( );
FILL FILL_0_AOI21X1_37 ( );
FILL FILL_1_AOI21X1_37 ( );
FILL FILL_2_AOI21X1_37 ( );
FILL FILL_3_AOI21X1_37 ( );
FILL FILL_4_AOI21X1_37 ( );
FILL FILL_5_AOI21X1_37 ( );
FILL FILL_6_AOI21X1_37 ( );
FILL FILL_7_AOI21X1_37 ( );
FILL FILL_8_AOI21X1_37 ( );
FILL FILL_9_AOI21X1_37 ( );
FILL FILL_0_OR2X2_3 ( );
FILL FILL_1_OR2X2_3 ( );
FILL FILL_2_OR2X2_3 ( );
FILL FILL_3_OR2X2_3 ( );
FILL FILL_4_OR2X2_3 ( );
FILL FILL_5_OR2X2_3 ( );
FILL FILL_6_OR2X2_3 ( );
FILL FILL_7_OR2X2_3 ( );
FILL FILL_8_OR2X2_3 ( );
FILL FILL_0_NAND3X1_229 ( );
FILL FILL_1_NAND3X1_229 ( );
FILL FILL_2_NAND3X1_229 ( );
FILL FILL_3_NAND3X1_229 ( );
FILL FILL_4_NAND3X1_229 ( );
FILL FILL_5_NAND3X1_229 ( );
FILL FILL_6_NAND3X1_229 ( );
FILL FILL_7_NAND3X1_229 ( );
FILL FILL_8_NAND3X1_229 ( );
FILL FILL_9_NAND3X1_229 ( );
FILL FILL_0_NAND3X1_228 ( );
FILL FILL_1_NAND3X1_228 ( );
FILL FILL_2_NAND3X1_228 ( );
FILL FILL_3_NAND3X1_228 ( );
FILL FILL_4_NAND3X1_228 ( );
FILL FILL_5_NAND3X1_228 ( );
FILL FILL_6_NAND3X1_228 ( );
FILL FILL_7_NAND3X1_228 ( );
FILL FILL_8_NAND3X1_228 ( );
FILL FILL_0_CLKBUF1_46 ( );
FILL FILL_1_CLKBUF1_46 ( );
FILL FILL_2_CLKBUF1_46 ( );
FILL FILL_3_CLKBUF1_46 ( );
FILL FILL_4_CLKBUF1_46 ( );
FILL FILL_5_CLKBUF1_46 ( );
FILL FILL_6_CLKBUF1_46 ( );
FILL FILL_7_CLKBUF1_46 ( );
FILL FILL_8_CLKBUF1_46 ( );
FILL FILL_9_CLKBUF1_46 ( );
FILL FILL_10_CLKBUF1_46 ( );
FILL FILL_11_CLKBUF1_46 ( );
FILL FILL_12_CLKBUF1_46 ( );
FILL FILL_13_CLKBUF1_46 ( );
FILL FILL_14_CLKBUF1_46 ( );
FILL FILL_15_CLKBUF1_46 ( );
FILL FILL_16_CLKBUF1_46 ( );
FILL FILL_17_CLKBUF1_46 ( );
FILL FILL_18_CLKBUF1_46 ( );
FILL FILL_19_CLKBUF1_46 ( );
FILL FILL_20_CLKBUF1_46 ( );
FILL FILL_0_DFFSR_52 ( );
FILL FILL_1_DFFSR_52 ( );
FILL FILL_2_DFFSR_52 ( );
FILL FILL_3_DFFSR_52 ( );
FILL FILL_4_DFFSR_52 ( );
FILL FILL_5_DFFSR_52 ( );
FILL FILL_6_DFFSR_52 ( );
FILL FILL_7_DFFSR_52 ( );
FILL FILL_8_DFFSR_52 ( );
FILL FILL_9_DFFSR_52 ( );
FILL FILL_10_DFFSR_52 ( );
FILL FILL_11_DFFSR_52 ( );
FILL FILL_12_DFFSR_52 ( );
FILL FILL_13_DFFSR_52 ( );
FILL FILL_14_DFFSR_52 ( );
FILL FILL_15_DFFSR_52 ( );
FILL FILL_16_DFFSR_52 ( );
FILL FILL_17_DFFSR_52 ( );
FILL FILL_18_DFFSR_52 ( );
FILL FILL_19_DFFSR_52 ( );
FILL FILL_20_DFFSR_52 ( );
FILL FILL_21_DFFSR_52 ( );
FILL FILL_22_DFFSR_52 ( );
FILL FILL_23_DFFSR_52 ( );
FILL FILL_24_DFFSR_52 ( );
FILL FILL_25_DFFSR_52 ( );
FILL FILL_26_DFFSR_52 ( );
FILL FILL_27_DFFSR_52 ( );
FILL FILL_28_DFFSR_52 ( );
FILL FILL_29_DFFSR_52 ( );
FILL FILL_30_DFFSR_52 ( );
FILL FILL_31_DFFSR_52 ( );
FILL FILL_32_DFFSR_52 ( );
FILL FILL_33_DFFSR_52 ( );
FILL FILL_34_DFFSR_52 ( );
FILL FILL_35_DFFSR_52 ( );
FILL FILL_36_DFFSR_52 ( );
FILL FILL_37_DFFSR_52 ( );
FILL FILL_38_DFFSR_52 ( );
FILL FILL_39_DFFSR_52 ( );
FILL FILL_40_DFFSR_52 ( );
FILL FILL_41_DFFSR_52 ( );
FILL FILL_42_DFFSR_52 ( );
FILL FILL_43_DFFSR_52 ( );
FILL FILL_44_DFFSR_52 ( );
FILL FILL_45_DFFSR_52 ( );
FILL FILL_46_DFFSR_52 ( );
FILL FILL_47_DFFSR_52 ( );
FILL FILL_48_DFFSR_52 ( );
FILL FILL_49_DFFSR_52 ( );
FILL FILL_50_DFFSR_52 ( );
FILL FILL_0_INVX1_11 ( );
FILL FILL_1_INVX1_11 ( );
FILL FILL_2_INVX1_11 ( );
FILL FILL_3_INVX1_11 ( );
FILL FILL_4_INVX1_11 ( );
FILL FILL_0_DFFSR_15 ( );
FILL FILL_1_DFFSR_15 ( );
FILL FILL_2_DFFSR_15 ( );
FILL FILL_3_DFFSR_15 ( );
FILL FILL_4_DFFSR_15 ( );
FILL FILL_5_DFFSR_15 ( );
FILL FILL_6_DFFSR_15 ( );
FILL FILL_7_DFFSR_15 ( );
FILL FILL_8_DFFSR_15 ( );
FILL FILL_9_DFFSR_15 ( );
FILL FILL_10_DFFSR_15 ( );
FILL FILL_11_DFFSR_15 ( );
FILL FILL_12_DFFSR_15 ( );
FILL FILL_13_DFFSR_15 ( );
FILL FILL_14_DFFSR_15 ( );
FILL FILL_15_DFFSR_15 ( );
FILL FILL_16_DFFSR_15 ( );
FILL FILL_17_DFFSR_15 ( );
FILL FILL_18_DFFSR_15 ( );
FILL FILL_19_DFFSR_15 ( );
FILL FILL_20_DFFSR_15 ( );
FILL FILL_21_DFFSR_15 ( );
FILL FILL_22_DFFSR_15 ( );
FILL FILL_23_DFFSR_15 ( );
FILL FILL_24_DFFSR_15 ( );
FILL FILL_25_DFFSR_15 ( );
FILL FILL_26_DFFSR_15 ( );
FILL FILL_27_DFFSR_15 ( );
FILL FILL_28_DFFSR_15 ( );
FILL FILL_29_DFFSR_15 ( );
FILL FILL_30_DFFSR_15 ( );
FILL FILL_31_DFFSR_15 ( );
FILL FILL_32_DFFSR_15 ( );
FILL FILL_33_DFFSR_15 ( );
FILL FILL_34_DFFSR_15 ( );
FILL FILL_35_DFFSR_15 ( );
FILL FILL_36_DFFSR_15 ( );
FILL FILL_37_DFFSR_15 ( );
FILL FILL_38_DFFSR_15 ( );
FILL FILL_39_DFFSR_15 ( );
FILL FILL_40_DFFSR_15 ( );
FILL FILL_41_DFFSR_15 ( );
FILL FILL_42_DFFSR_15 ( );
FILL FILL_43_DFFSR_15 ( );
FILL FILL_44_DFFSR_15 ( );
FILL FILL_45_DFFSR_15 ( );
FILL FILL_46_DFFSR_15 ( );
FILL FILL_47_DFFSR_15 ( );
FILL FILL_48_DFFSR_15 ( );
FILL FILL_49_DFFSR_15 ( );
FILL FILL_50_DFFSR_15 ( );
FILL FILL_0_INVX1_45 ( );
FILL FILL_1_INVX1_45 ( );
FILL FILL_2_INVX1_45 ( );
FILL FILL_3_INVX1_45 ( );
FILL FILL_0_OAI22X1_4 ( );
FILL FILL_1_OAI22X1_4 ( );
FILL FILL_2_OAI22X1_4 ( );
FILL FILL_3_OAI22X1_4 ( );
FILL FILL_4_OAI22X1_4 ( );
FILL FILL_5_OAI22X1_4 ( );
FILL FILL_6_OAI22X1_4 ( );
FILL FILL_7_OAI22X1_4 ( );
FILL FILL_8_OAI22X1_4 ( );
FILL FILL_9_OAI22X1_4 ( );
FILL FILL_10_OAI22X1_4 ( );
FILL FILL_11_OAI22X1_4 ( );
FILL FILL_0_NAND2X1_24 ( );
FILL FILL_1_NAND2X1_24 ( );
FILL FILL_2_NAND2X1_24 ( );
FILL FILL_3_NAND2X1_24 ( );
FILL FILL_4_NAND2X1_24 ( );
FILL FILL_5_NAND2X1_24 ( );
FILL FILL_6_NAND2X1_24 ( );
FILL FILL_0_DFFSR_78 ( );
FILL FILL_1_DFFSR_78 ( );
FILL FILL_2_DFFSR_78 ( );
FILL FILL_3_DFFSR_78 ( );
FILL FILL_4_DFFSR_78 ( );
FILL FILL_5_DFFSR_78 ( );
FILL FILL_6_DFFSR_78 ( );
FILL FILL_7_DFFSR_78 ( );
FILL FILL_8_DFFSR_78 ( );
FILL FILL_9_DFFSR_78 ( );
FILL FILL_10_DFFSR_78 ( );
FILL FILL_11_DFFSR_78 ( );
FILL FILL_12_DFFSR_78 ( );
FILL FILL_13_DFFSR_78 ( );
FILL FILL_14_DFFSR_78 ( );
FILL FILL_15_DFFSR_78 ( );
FILL FILL_16_DFFSR_78 ( );
FILL FILL_17_DFFSR_78 ( );
FILL FILL_18_DFFSR_78 ( );
FILL FILL_19_DFFSR_78 ( );
FILL FILL_20_DFFSR_78 ( );
FILL FILL_21_DFFSR_78 ( );
FILL FILL_22_DFFSR_78 ( );
FILL FILL_23_DFFSR_78 ( );
FILL FILL_24_DFFSR_78 ( );
FILL FILL_25_DFFSR_78 ( );
FILL FILL_26_DFFSR_78 ( );
FILL FILL_27_DFFSR_78 ( );
FILL FILL_28_DFFSR_78 ( );
FILL FILL_29_DFFSR_78 ( );
FILL FILL_30_DFFSR_78 ( );
FILL FILL_31_DFFSR_78 ( );
FILL FILL_32_DFFSR_78 ( );
FILL FILL_33_DFFSR_78 ( );
FILL FILL_34_DFFSR_78 ( );
FILL FILL_35_DFFSR_78 ( );
FILL FILL_36_DFFSR_78 ( );
FILL FILL_37_DFFSR_78 ( );
FILL FILL_38_DFFSR_78 ( );
FILL FILL_39_DFFSR_78 ( );
FILL FILL_40_DFFSR_78 ( );
FILL FILL_41_DFFSR_78 ( );
FILL FILL_42_DFFSR_78 ( );
FILL FILL_43_DFFSR_78 ( );
FILL FILL_44_DFFSR_78 ( );
FILL FILL_45_DFFSR_78 ( );
FILL FILL_46_DFFSR_78 ( );
FILL FILL_47_DFFSR_78 ( );
FILL FILL_48_DFFSR_78 ( );
FILL FILL_49_DFFSR_78 ( );
FILL FILL_50_DFFSR_78 ( );
FILL FILL_51_DFFSR_78 ( );
FILL FILL_0_NAND3X1_47 ( );
FILL FILL_1_NAND3X1_47 ( );
FILL FILL_2_NAND3X1_47 ( );
FILL FILL_3_NAND3X1_47 ( );
FILL FILL_4_NAND3X1_47 ( );
FILL FILL_5_NAND3X1_47 ( );
FILL FILL_6_NAND3X1_47 ( );
FILL FILL_7_NAND3X1_47 ( );
FILL FILL_8_NAND3X1_47 ( );
FILL FILL_0_DFFPOSX1_7 ( );
FILL FILL_1_DFFPOSX1_7 ( );
FILL FILL_2_DFFPOSX1_7 ( );
FILL FILL_3_DFFPOSX1_7 ( );
FILL FILL_4_DFFPOSX1_7 ( );
FILL FILL_5_DFFPOSX1_7 ( );
FILL FILL_6_DFFPOSX1_7 ( );
FILL FILL_7_DFFPOSX1_7 ( );
FILL FILL_8_DFFPOSX1_7 ( );
FILL FILL_9_DFFPOSX1_7 ( );
FILL FILL_10_DFFPOSX1_7 ( );
FILL FILL_11_DFFPOSX1_7 ( );
FILL FILL_12_DFFPOSX1_7 ( );
FILL FILL_13_DFFPOSX1_7 ( );
FILL FILL_14_DFFPOSX1_7 ( );
FILL FILL_15_DFFPOSX1_7 ( );
FILL FILL_16_DFFPOSX1_7 ( );
FILL FILL_17_DFFPOSX1_7 ( );
FILL FILL_18_DFFPOSX1_7 ( );
FILL FILL_19_DFFPOSX1_7 ( );
FILL FILL_20_DFFPOSX1_7 ( );
FILL FILL_21_DFFPOSX1_7 ( );
FILL FILL_22_DFFPOSX1_7 ( );
FILL FILL_23_DFFPOSX1_7 ( );
FILL FILL_24_DFFPOSX1_7 ( );
FILL FILL_25_DFFPOSX1_7 ( );
FILL FILL_26_DFFPOSX1_7 ( );
FILL FILL_27_DFFPOSX1_7 ( );
FILL FILL_0_DFFSR_110 ( );
FILL FILL_1_DFFSR_110 ( );
FILL FILL_2_DFFSR_110 ( );
FILL FILL_3_DFFSR_110 ( );
FILL FILL_4_DFFSR_110 ( );
FILL FILL_5_DFFSR_110 ( );
FILL FILL_6_DFFSR_110 ( );
FILL FILL_7_DFFSR_110 ( );
FILL FILL_8_DFFSR_110 ( );
FILL FILL_9_DFFSR_110 ( );
FILL FILL_10_DFFSR_110 ( );
FILL FILL_11_DFFSR_110 ( );
FILL FILL_12_DFFSR_110 ( );
FILL FILL_13_DFFSR_110 ( );
FILL FILL_14_DFFSR_110 ( );
FILL FILL_15_DFFSR_110 ( );
FILL FILL_16_DFFSR_110 ( );
FILL FILL_17_DFFSR_110 ( );
FILL FILL_18_DFFSR_110 ( );
FILL FILL_19_DFFSR_110 ( );
FILL FILL_20_DFFSR_110 ( );
FILL FILL_21_DFFSR_110 ( );
FILL FILL_22_DFFSR_110 ( );
FILL FILL_23_DFFSR_110 ( );
FILL FILL_24_DFFSR_110 ( );
FILL FILL_25_DFFSR_110 ( );
FILL FILL_26_DFFSR_110 ( );
FILL FILL_27_DFFSR_110 ( );
FILL FILL_28_DFFSR_110 ( );
FILL FILL_29_DFFSR_110 ( );
FILL FILL_30_DFFSR_110 ( );
FILL FILL_31_DFFSR_110 ( );
FILL FILL_32_DFFSR_110 ( );
FILL FILL_33_DFFSR_110 ( );
FILL FILL_34_DFFSR_110 ( );
FILL FILL_35_DFFSR_110 ( );
FILL FILL_36_DFFSR_110 ( );
FILL FILL_37_DFFSR_110 ( );
FILL FILL_38_DFFSR_110 ( );
FILL FILL_39_DFFSR_110 ( );
FILL FILL_40_DFFSR_110 ( );
FILL FILL_41_DFFSR_110 ( );
FILL FILL_42_DFFSR_110 ( );
FILL FILL_43_DFFSR_110 ( );
FILL FILL_44_DFFSR_110 ( );
FILL FILL_45_DFFSR_110 ( );
FILL FILL_46_DFFSR_110 ( );
FILL FILL_47_DFFSR_110 ( );
FILL FILL_48_DFFSR_110 ( );
FILL FILL_49_DFFSR_110 ( );
FILL FILL_50_DFFSR_110 ( );
FILL FILL_0_INVX1_36 ( );
FILL FILL_1_INVX1_36 ( );
FILL FILL_2_INVX1_36 ( );
FILL FILL_3_INVX1_36 ( );
FILL FILL_4_INVX1_36 ( );
FILL FILL_0_BUFX2_51 ( );
FILL FILL_1_BUFX2_51 ( );
FILL FILL_2_BUFX2_51 ( );
FILL FILL_3_BUFX2_51 ( );
FILL FILL_4_BUFX2_51 ( );
FILL FILL_5_BUFX2_51 ( );
FILL FILL_6_BUFX2_51 ( );
FILL FILL_0_CLKBUF1_16 ( );
FILL FILL_1_CLKBUF1_16 ( );
FILL FILL_2_CLKBUF1_16 ( );
FILL FILL_3_CLKBUF1_16 ( );
FILL FILL_4_CLKBUF1_16 ( );
FILL FILL_5_CLKBUF1_16 ( );
FILL FILL_6_CLKBUF1_16 ( );
FILL FILL_7_CLKBUF1_16 ( );
FILL FILL_8_CLKBUF1_16 ( );
FILL FILL_9_CLKBUF1_16 ( );
FILL FILL_10_CLKBUF1_16 ( );
FILL FILL_11_CLKBUF1_16 ( );
FILL FILL_12_CLKBUF1_16 ( );
FILL FILL_13_CLKBUF1_16 ( );
FILL FILL_14_CLKBUF1_16 ( );
FILL FILL_15_CLKBUF1_16 ( );
FILL FILL_16_CLKBUF1_16 ( );
FILL FILL_17_CLKBUF1_16 ( );
FILL FILL_18_CLKBUF1_16 ( );
FILL FILL_19_CLKBUF1_16 ( );
FILL FILL_20_CLKBUF1_16 ( );
FILL FILL_0_DFFSR_101 ( );
FILL FILL_1_DFFSR_101 ( );
FILL FILL_2_DFFSR_101 ( );
FILL FILL_3_DFFSR_101 ( );
FILL FILL_4_DFFSR_101 ( );
FILL FILL_5_DFFSR_101 ( );
FILL FILL_6_DFFSR_101 ( );
FILL FILL_7_DFFSR_101 ( );
FILL FILL_8_DFFSR_101 ( );
FILL FILL_9_DFFSR_101 ( );
FILL FILL_10_DFFSR_101 ( );
FILL FILL_11_DFFSR_101 ( );
FILL FILL_12_DFFSR_101 ( );
FILL FILL_13_DFFSR_101 ( );
FILL FILL_14_DFFSR_101 ( );
FILL FILL_15_DFFSR_101 ( );
FILL FILL_16_DFFSR_101 ( );
FILL FILL_17_DFFSR_101 ( );
FILL FILL_18_DFFSR_101 ( );
FILL FILL_19_DFFSR_101 ( );
FILL FILL_20_DFFSR_101 ( );
FILL FILL_21_DFFSR_101 ( );
FILL FILL_22_DFFSR_101 ( );
FILL FILL_23_DFFSR_101 ( );
FILL FILL_24_DFFSR_101 ( );
FILL FILL_25_DFFSR_101 ( );
FILL FILL_26_DFFSR_101 ( );
FILL FILL_27_DFFSR_101 ( );
FILL FILL_28_DFFSR_101 ( );
FILL FILL_29_DFFSR_101 ( );
FILL FILL_30_DFFSR_101 ( );
FILL FILL_31_DFFSR_101 ( );
FILL FILL_32_DFFSR_101 ( );
FILL FILL_33_DFFSR_101 ( );
FILL FILL_34_DFFSR_101 ( );
FILL FILL_35_DFFSR_101 ( );
FILL FILL_36_DFFSR_101 ( );
FILL FILL_37_DFFSR_101 ( );
FILL FILL_38_DFFSR_101 ( );
FILL FILL_39_DFFSR_101 ( );
FILL FILL_40_DFFSR_101 ( );
FILL FILL_41_DFFSR_101 ( );
FILL FILL_42_DFFSR_101 ( );
FILL FILL_43_DFFSR_101 ( );
FILL FILL_44_DFFSR_101 ( );
FILL FILL_45_DFFSR_101 ( );
FILL FILL_46_DFFSR_101 ( );
FILL FILL_47_DFFSR_101 ( );
FILL FILL_48_DFFSR_101 ( );
FILL FILL_49_DFFSR_101 ( );
FILL FILL_50_DFFSR_101 ( );
FILL FILL_51_DFFSR_101 ( );
FILL FILL_0_DFFSR_234 ( );
FILL FILL_1_DFFSR_234 ( );
FILL FILL_2_DFFSR_234 ( );
FILL FILL_3_DFFSR_234 ( );
FILL FILL_4_DFFSR_234 ( );
FILL FILL_5_DFFSR_234 ( );
FILL FILL_6_DFFSR_234 ( );
FILL FILL_7_DFFSR_234 ( );
FILL FILL_8_DFFSR_234 ( );
FILL FILL_9_DFFSR_234 ( );
FILL FILL_10_DFFSR_234 ( );
FILL FILL_11_DFFSR_234 ( );
FILL FILL_12_DFFSR_234 ( );
FILL FILL_13_DFFSR_234 ( );
FILL FILL_14_DFFSR_234 ( );
FILL FILL_15_DFFSR_234 ( );
FILL FILL_16_DFFSR_234 ( );
FILL FILL_17_DFFSR_234 ( );
FILL FILL_18_DFFSR_234 ( );
FILL FILL_19_DFFSR_234 ( );
FILL FILL_20_DFFSR_234 ( );
FILL FILL_21_DFFSR_234 ( );
FILL FILL_22_DFFSR_234 ( );
FILL FILL_23_DFFSR_234 ( );
FILL FILL_24_DFFSR_234 ( );
FILL FILL_25_DFFSR_234 ( );
FILL FILL_26_DFFSR_234 ( );
FILL FILL_27_DFFSR_234 ( );
FILL FILL_28_DFFSR_234 ( );
FILL FILL_29_DFFSR_234 ( );
FILL FILL_30_DFFSR_234 ( );
FILL FILL_31_DFFSR_234 ( );
FILL FILL_32_DFFSR_234 ( );
FILL FILL_33_DFFSR_234 ( );
FILL FILL_34_DFFSR_234 ( );
FILL FILL_35_DFFSR_234 ( );
FILL FILL_36_DFFSR_234 ( );
FILL FILL_37_DFFSR_234 ( );
FILL FILL_38_DFFSR_234 ( );
FILL FILL_39_DFFSR_234 ( );
FILL FILL_40_DFFSR_234 ( );
FILL FILL_41_DFFSR_234 ( );
FILL FILL_42_DFFSR_234 ( );
FILL FILL_43_DFFSR_234 ( );
FILL FILL_44_DFFSR_234 ( );
FILL FILL_45_DFFSR_234 ( );
FILL FILL_46_DFFSR_234 ( );
FILL FILL_47_DFFSR_234 ( );
FILL FILL_48_DFFSR_234 ( );
FILL FILL_49_DFFSR_234 ( );
FILL FILL_50_DFFSR_234 ( );
FILL FILL_0_NAND3X1_235 ( );
FILL FILL_1_NAND3X1_235 ( );
FILL FILL_2_NAND3X1_235 ( );
FILL FILL_3_NAND3X1_235 ( );
FILL FILL_4_NAND3X1_235 ( );
FILL FILL_5_NAND3X1_235 ( );
FILL FILL_6_NAND3X1_235 ( );
FILL FILL_7_NAND3X1_235 ( );
FILL FILL_8_NAND3X1_235 ( );
FILL FILL_0_NAND3X1_227 ( );
FILL FILL_1_NAND3X1_227 ( );
FILL FILL_2_NAND3X1_227 ( );
FILL FILL_3_NAND3X1_227 ( );
FILL FILL_4_NAND3X1_227 ( );
FILL FILL_5_NAND3X1_227 ( );
FILL FILL_6_NAND3X1_227 ( );
FILL FILL_7_NAND3X1_227 ( );
FILL FILL_8_NAND3X1_227 ( );
FILL FILL_0_NAND3X1_233 ( );
FILL FILL_1_NAND3X1_233 ( );
FILL FILL_2_NAND3X1_233 ( );
FILL FILL_3_NAND3X1_233 ( );
FILL FILL_4_NAND3X1_233 ( );
FILL FILL_5_NAND3X1_233 ( );
FILL FILL_6_NAND3X1_233 ( );
FILL FILL_7_NAND3X1_233 ( );
FILL FILL_8_NAND3X1_233 ( );
FILL FILL_0_NAND3X1_230 ( );
FILL FILL_1_NAND3X1_230 ( );
FILL FILL_2_NAND3X1_230 ( );
FILL FILL_3_NAND3X1_230 ( );
FILL FILL_4_NAND3X1_230 ( );
FILL FILL_5_NAND3X1_230 ( );
FILL FILL_6_NAND3X1_230 ( );
FILL FILL_7_NAND3X1_230 ( );
FILL FILL_8_NAND3X1_230 ( );
FILL FILL_0_NAND3X1_225 ( );
FILL FILL_1_NAND3X1_225 ( );
FILL FILL_2_NAND3X1_225 ( );
FILL FILL_3_NAND3X1_225 ( );
FILL FILL_4_NAND3X1_225 ( );
FILL FILL_5_NAND3X1_225 ( );
FILL FILL_6_NAND3X1_225 ( );
FILL FILL_7_NAND3X1_225 ( );
FILL FILL_8_NAND3X1_225 ( );
FILL FILL_9_NAND3X1_225 ( );
FILL FILL_0_DFFSR_4 ( );
FILL FILL_1_DFFSR_4 ( );
FILL FILL_2_DFFSR_4 ( );
FILL FILL_3_DFFSR_4 ( );
FILL FILL_4_DFFSR_4 ( );
FILL FILL_5_DFFSR_4 ( );
FILL FILL_6_DFFSR_4 ( );
FILL FILL_7_DFFSR_4 ( );
FILL FILL_8_DFFSR_4 ( );
FILL FILL_9_DFFSR_4 ( );
FILL FILL_10_DFFSR_4 ( );
FILL FILL_11_DFFSR_4 ( );
FILL FILL_12_DFFSR_4 ( );
FILL FILL_13_DFFSR_4 ( );
FILL FILL_14_DFFSR_4 ( );
FILL FILL_15_DFFSR_4 ( );
FILL FILL_16_DFFSR_4 ( );
FILL FILL_17_DFFSR_4 ( );
FILL FILL_18_DFFSR_4 ( );
FILL FILL_19_DFFSR_4 ( );
FILL FILL_20_DFFSR_4 ( );
FILL FILL_21_DFFSR_4 ( );
FILL FILL_22_DFFSR_4 ( );
FILL FILL_23_DFFSR_4 ( );
FILL FILL_24_DFFSR_4 ( );
FILL FILL_25_DFFSR_4 ( );
FILL FILL_26_DFFSR_4 ( );
FILL FILL_27_DFFSR_4 ( );
FILL FILL_28_DFFSR_4 ( );
FILL FILL_29_DFFSR_4 ( );
FILL FILL_30_DFFSR_4 ( );
FILL FILL_31_DFFSR_4 ( );
FILL FILL_32_DFFSR_4 ( );
FILL FILL_33_DFFSR_4 ( );
FILL FILL_34_DFFSR_4 ( );
FILL FILL_35_DFFSR_4 ( );
FILL FILL_36_DFFSR_4 ( );
FILL FILL_37_DFFSR_4 ( );
FILL FILL_38_DFFSR_4 ( );
FILL FILL_39_DFFSR_4 ( );
FILL FILL_40_DFFSR_4 ( );
FILL FILL_41_DFFSR_4 ( );
FILL FILL_42_DFFSR_4 ( );
FILL FILL_43_DFFSR_4 ( );
FILL FILL_44_DFFSR_4 ( );
FILL FILL_45_DFFSR_4 ( );
FILL FILL_46_DFFSR_4 ( );
FILL FILL_47_DFFSR_4 ( );
FILL FILL_48_DFFSR_4 ( );
FILL FILL_49_DFFSR_4 ( );
FILL FILL_50_DFFSR_4 ( );
FILL FILL_0_BUFX2_78 ( );
FILL FILL_1_BUFX2_78 ( );
FILL FILL_2_BUFX2_78 ( );
FILL FILL_3_BUFX2_78 ( );
FILL FILL_4_BUFX2_78 ( );
FILL FILL_5_BUFX2_78 ( );
FILL FILL_6_BUFX2_78 ( );
FILL FILL_0_DFFPOSX1_11 ( );
FILL FILL_1_DFFPOSX1_11 ( );
FILL FILL_2_DFFPOSX1_11 ( );
FILL FILL_3_DFFPOSX1_11 ( );
FILL FILL_4_DFFPOSX1_11 ( );
FILL FILL_5_DFFPOSX1_11 ( );
FILL FILL_6_DFFPOSX1_11 ( );
FILL FILL_7_DFFPOSX1_11 ( );
FILL FILL_8_DFFPOSX1_11 ( );
FILL FILL_9_DFFPOSX1_11 ( );
FILL FILL_10_DFFPOSX1_11 ( );
FILL FILL_11_DFFPOSX1_11 ( );
FILL FILL_12_DFFPOSX1_11 ( );
FILL FILL_13_DFFPOSX1_11 ( );
FILL FILL_14_DFFPOSX1_11 ( );
FILL FILL_15_DFFPOSX1_11 ( );
FILL FILL_16_DFFPOSX1_11 ( );
FILL FILL_17_DFFPOSX1_11 ( );
FILL FILL_18_DFFPOSX1_11 ( );
FILL FILL_19_DFFPOSX1_11 ( );
FILL FILL_20_DFFPOSX1_11 ( );
FILL FILL_21_DFFPOSX1_11 ( );
FILL FILL_22_DFFPOSX1_11 ( );
FILL FILL_23_DFFPOSX1_11 ( );
FILL FILL_24_DFFPOSX1_11 ( );
FILL FILL_25_DFFPOSX1_11 ( );
FILL FILL_26_DFFPOSX1_11 ( );
FILL FILL_27_DFFPOSX1_11 ( );
FILL FILL_0_DFFSR_55 ( );
FILL FILL_1_DFFSR_55 ( );
FILL FILL_2_DFFSR_55 ( );
FILL FILL_3_DFFSR_55 ( );
FILL FILL_4_DFFSR_55 ( );
FILL FILL_5_DFFSR_55 ( );
FILL FILL_6_DFFSR_55 ( );
FILL FILL_7_DFFSR_55 ( );
FILL FILL_8_DFFSR_55 ( );
FILL FILL_9_DFFSR_55 ( );
FILL FILL_10_DFFSR_55 ( );
FILL FILL_11_DFFSR_55 ( );
FILL FILL_12_DFFSR_55 ( );
FILL FILL_13_DFFSR_55 ( );
FILL FILL_14_DFFSR_55 ( );
FILL FILL_15_DFFSR_55 ( );
FILL FILL_16_DFFSR_55 ( );
FILL FILL_17_DFFSR_55 ( );
FILL FILL_18_DFFSR_55 ( );
FILL FILL_19_DFFSR_55 ( );
FILL FILL_20_DFFSR_55 ( );
FILL FILL_21_DFFSR_55 ( );
FILL FILL_22_DFFSR_55 ( );
FILL FILL_23_DFFSR_55 ( );
FILL FILL_24_DFFSR_55 ( );
FILL FILL_25_DFFSR_55 ( );
FILL FILL_26_DFFSR_55 ( );
FILL FILL_27_DFFSR_55 ( );
FILL FILL_28_DFFSR_55 ( );
FILL FILL_29_DFFSR_55 ( );
FILL FILL_30_DFFSR_55 ( );
FILL FILL_31_DFFSR_55 ( );
FILL FILL_32_DFFSR_55 ( );
FILL FILL_33_DFFSR_55 ( );
FILL FILL_34_DFFSR_55 ( );
FILL FILL_35_DFFSR_55 ( );
FILL FILL_36_DFFSR_55 ( );
FILL FILL_37_DFFSR_55 ( );
FILL FILL_38_DFFSR_55 ( );
FILL FILL_39_DFFSR_55 ( );
FILL FILL_40_DFFSR_55 ( );
FILL FILL_41_DFFSR_55 ( );
FILL FILL_42_DFFSR_55 ( );
FILL FILL_43_DFFSR_55 ( );
FILL FILL_44_DFFSR_55 ( );
FILL FILL_45_DFFSR_55 ( );
FILL FILL_46_DFFSR_55 ( );
FILL FILL_47_DFFSR_55 ( );
FILL FILL_48_DFFSR_55 ( );
FILL FILL_49_DFFSR_55 ( );
FILL FILL_50_DFFSR_55 ( );
FILL FILL_0_INVX1_46 ( );
FILL FILL_1_INVX1_46 ( );
FILL FILL_2_INVX1_46 ( );
FILL FILL_3_INVX1_46 ( );
FILL FILL_4_INVX1_46 ( );
FILL FILL_0_NOR2X1_24 ( );
FILL FILL_1_NOR2X1_24 ( );
FILL FILL_2_NOR2X1_24 ( );
FILL FILL_3_NOR2X1_24 ( );
FILL FILL_4_NOR2X1_24 ( );
FILL FILL_5_NOR2X1_24 ( );
FILL FILL_6_NOR2X1_24 ( );
FILL FILL_0_NOR2X1_9 ( );
FILL FILL_1_NOR2X1_9 ( );
FILL FILL_2_NOR2X1_9 ( );
FILL FILL_3_NOR2X1_9 ( );
FILL FILL_4_NOR2X1_9 ( );
FILL FILL_5_NOR2X1_9 ( );
FILL FILL_6_NOR2X1_9 ( );
FILL FILL_0_DFFSR_86 ( );
FILL FILL_1_DFFSR_86 ( );
FILL FILL_2_DFFSR_86 ( );
FILL FILL_3_DFFSR_86 ( );
FILL FILL_4_DFFSR_86 ( );
FILL FILL_5_DFFSR_86 ( );
FILL FILL_6_DFFSR_86 ( );
FILL FILL_7_DFFSR_86 ( );
FILL FILL_8_DFFSR_86 ( );
FILL FILL_9_DFFSR_86 ( );
FILL FILL_10_DFFSR_86 ( );
FILL FILL_11_DFFSR_86 ( );
FILL FILL_12_DFFSR_86 ( );
FILL FILL_13_DFFSR_86 ( );
FILL FILL_14_DFFSR_86 ( );
FILL FILL_15_DFFSR_86 ( );
FILL FILL_16_DFFSR_86 ( );
FILL FILL_17_DFFSR_86 ( );
FILL FILL_18_DFFSR_86 ( );
FILL FILL_19_DFFSR_86 ( );
FILL FILL_20_DFFSR_86 ( );
FILL FILL_21_DFFSR_86 ( );
FILL FILL_22_DFFSR_86 ( );
FILL FILL_23_DFFSR_86 ( );
FILL FILL_24_DFFSR_86 ( );
FILL FILL_25_DFFSR_86 ( );
FILL FILL_26_DFFSR_86 ( );
FILL FILL_27_DFFSR_86 ( );
FILL FILL_28_DFFSR_86 ( );
FILL FILL_29_DFFSR_86 ( );
FILL FILL_30_DFFSR_86 ( );
FILL FILL_31_DFFSR_86 ( );
FILL FILL_32_DFFSR_86 ( );
FILL FILL_33_DFFSR_86 ( );
FILL FILL_34_DFFSR_86 ( );
FILL FILL_35_DFFSR_86 ( );
FILL FILL_36_DFFSR_86 ( );
FILL FILL_37_DFFSR_86 ( );
FILL FILL_38_DFFSR_86 ( );
FILL FILL_39_DFFSR_86 ( );
FILL FILL_40_DFFSR_86 ( );
FILL FILL_41_DFFSR_86 ( );
FILL FILL_42_DFFSR_86 ( );
FILL FILL_43_DFFSR_86 ( );
FILL FILL_44_DFFSR_86 ( );
FILL FILL_45_DFFSR_86 ( );
FILL FILL_46_DFFSR_86 ( );
FILL FILL_47_DFFSR_86 ( );
FILL FILL_48_DFFSR_86 ( );
FILL FILL_49_DFFSR_86 ( );
FILL FILL_50_DFFSR_86 ( );
FILL FILL_51_DFFSR_86 ( );
FILL FILL_0_NAND3X1_46 ( );
FILL FILL_1_NAND3X1_46 ( );
FILL FILL_2_NAND3X1_46 ( );
FILL FILL_3_NAND3X1_46 ( );
FILL FILL_4_NAND3X1_46 ( );
FILL FILL_5_NAND3X1_46 ( );
FILL FILL_6_NAND3X1_46 ( );
FILL FILL_7_NAND3X1_46 ( );
FILL FILL_8_NAND3X1_46 ( );
FILL FILL_0_NAND3X1_13 ( );
FILL FILL_1_NAND3X1_13 ( );
FILL FILL_2_NAND3X1_13 ( );
FILL FILL_3_NAND3X1_13 ( );
FILL FILL_4_NAND3X1_13 ( );
FILL FILL_5_NAND3X1_13 ( );
FILL FILL_6_NAND3X1_13 ( );
FILL FILL_7_NAND3X1_13 ( );
FILL FILL_8_NAND3X1_13 ( );
FILL FILL_9_NAND3X1_13 ( );
FILL FILL_0_AOI22X1_6 ( );
FILL FILL_1_AOI22X1_6 ( );
FILL FILL_2_AOI22X1_6 ( );
FILL FILL_3_AOI22X1_6 ( );
FILL FILL_4_AOI22X1_6 ( );
FILL FILL_5_AOI22X1_6 ( );
FILL FILL_6_AOI22X1_6 ( );
FILL FILL_7_AOI22X1_6 ( );
FILL FILL_8_AOI22X1_6 ( );
FILL FILL_9_AOI22X1_6 ( );
FILL FILL_10_AOI22X1_6 ( );
FILL FILL_11_AOI22X1_6 ( );
FILL FILL_0_NAND3X1_14 ( );
FILL FILL_1_NAND3X1_14 ( );
FILL FILL_2_NAND3X1_14 ( );
FILL FILL_3_NAND3X1_14 ( );
FILL FILL_4_NAND3X1_14 ( );
FILL FILL_5_NAND3X1_14 ( );
FILL FILL_6_NAND3X1_14 ( );
FILL FILL_7_NAND3X1_14 ( );
FILL FILL_8_NAND3X1_14 ( );
FILL FILL_0_NAND3X1_15 ( );
FILL FILL_1_NAND3X1_15 ( );
FILL FILL_2_NAND3X1_15 ( );
FILL FILL_3_NAND3X1_15 ( );
FILL FILL_4_NAND3X1_15 ( );
FILL FILL_5_NAND3X1_15 ( );
FILL FILL_6_NAND3X1_15 ( );
FILL FILL_7_NAND3X1_15 ( );
FILL FILL_8_NAND3X1_15 ( );
FILL FILL_0_OAI22X1_23 ( );
FILL FILL_1_OAI22X1_23 ( );
FILL FILL_2_OAI22X1_23 ( );
FILL FILL_3_OAI22X1_23 ( );
FILL FILL_4_OAI22X1_23 ( );
FILL FILL_5_OAI22X1_23 ( );
FILL FILL_6_OAI22X1_23 ( );
FILL FILL_7_OAI22X1_23 ( );
FILL FILL_8_OAI22X1_23 ( );
FILL FILL_9_OAI22X1_23 ( );
FILL FILL_10_OAI22X1_23 ( );
FILL FILL_0_DFFSR_80 ( );
FILL FILL_1_DFFSR_80 ( );
FILL FILL_2_DFFSR_80 ( );
FILL FILL_3_DFFSR_80 ( );
FILL FILL_4_DFFSR_80 ( );
FILL FILL_5_DFFSR_80 ( );
FILL FILL_6_DFFSR_80 ( );
FILL FILL_7_DFFSR_80 ( );
FILL FILL_8_DFFSR_80 ( );
FILL FILL_9_DFFSR_80 ( );
FILL FILL_10_DFFSR_80 ( );
FILL FILL_11_DFFSR_80 ( );
FILL FILL_12_DFFSR_80 ( );
FILL FILL_13_DFFSR_80 ( );
FILL FILL_14_DFFSR_80 ( );
FILL FILL_15_DFFSR_80 ( );
FILL FILL_16_DFFSR_80 ( );
FILL FILL_17_DFFSR_80 ( );
FILL FILL_18_DFFSR_80 ( );
FILL FILL_19_DFFSR_80 ( );
FILL FILL_20_DFFSR_80 ( );
FILL FILL_21_DFFSR_80 ( );
FILL FILL_22_DFFSR_80 ( );
FILL FILL_23_DFFSR_80 ( );
FILL FILL_24_DFFSR_80 ( );
FILL FILL_25_DFFSR_80 ( );
FILL FILL_26_DFFSR_80 ( );
FILL FILL_27_DFFSR_80 ( );
FILL FILL_28_DFFSR_80 ( );
FILL FILL_29_DFFSR_80 ( );
FILL FILL_30_DFFSR_80 ( );
FILL FILL_31_DFFSR_80 ( );
FILL FILL_32_DFFSR_80 ( );
FILL FILL_33_DFFSR_80 ( );
FILL FILL_34_DFFSR_80 ( );
FILL FILL_35_DFFSR_80 ( );
FILL FILL_36_DFFSR_80 ( );
FILL FILL_37_DFFSR_80 ( );
FILL FILL_38_DFFSR_80 ( );
FILL FILL_39_DFFSR_80 ( );
FILL FILL_40_DFFSR_80 ( );
FILL FILL_41_DFFSR_80 ( );
FILL FILL_42_DFFSR_80 ( );
FILL FILL_43_DFFSR_80 ( );
FILL FILL_44_DFFSR_80 ( );
FILL FILL_45_DFFSR_80 ( );
FILL FILL_46_DFFSR_80 ( );
FILL FILL_47_DFFSR_80 ( );
FILL FILL_48_DFFSR_80 ( );
FILL FILL_49_DFFSR_80 ( );
FILL FILL_50_DFFSR_80 ( );
FILL FILL_0_INVX1_54 ( );
FILL FILL_1_INVX1_54 ( );
FILL FILL_2_INVX1_54 ( );
FILL FILL_3_INVX1_54 ( );
FILL FILL_4_INVX1_54 ( );
FILL FILL_0_DFFSR_109 ( );
FILL FILL_1_DFFSR_109 ( );
FILL FILL_2_DFFSR_109 ( );
FILL FILL_3_DFFSR_109 ( );
FILL FILL_4_DFFSR_109 ( );
FILL FILL_5_DFFSR_109 ( );
FILL FILL_6_DFFSR_109 ( );
FILL FILL_7_DFFSR_109 ( );
FILL FILL_8_DFFSR_109 ( );
FILL FILL_9_DFFSR_109 ( );
FILL FILL_10_DFFSR_109 ( );
FILL FILL_11_DFFSR_109 ( );
FILL FILL_12_DFFSR_109 ( );
FILL FILL_13_DFFSR_109 ( );
FILL FILL_14_DFFSR_109 ( );
FILL FILL_15_DFFSR_109 ( );
FILL FILL_16_DFFSR_109 ( );
FILL FILL_17_DFFSR_109 ( );
FILL FILL_18_DFFSR_109 ( );
FILL FILL_19_DFFSR_109 ( );
FILL FILL_20_DFFSR_109 ( );
FILL FILL_21_DFFSR_109 ( );
FILL FILL_22_DFFSR_109 ( );
FILL FILL_23_DFFSR_109 ( );
FILL FILL_24_DFFSR_109 ( );
FILL FILL_25_DFFSR_109 ( );
FILL FILL_26_DFFSR_109 ( );
FILL FILL_27_DFFSR_109 ( );
FILL FILL_28_DFFSR_109 ( );
FILL FILL_29_DFFSR_109 ( );
FILL FILL_30_DFFSR_109 ( );
FILL FILL_31_DFFSR_109 ( );
FILL FILL_32_DFFSR_109 ( );
FILL FILL_33_DFFSR_109 ( );
FILL FILL_34_DFFSR_109 ( );
FILL FILL_35_DFFSR_109 ( );
FILL FILL_36_DFFSR_109 ( );
FILL FILL_37_DFFSR_109 ( );
FILL FILL_38_DFFSR_109 ( );
FILL FILL_39_DFFSR_109 ( );
FILL FILL_40_DFFSR_109 ( );
FILL FILL_41_DFFSR_109 ( );
FILL FILL_42_DFFSR_109 ( );
FILL FILL_43_DFFSR_109 ( );
FILL FILL_44_DFFSR_109 ( );
FILL FILL_45_DFFSR_109 ( );
FILL FILL_46_DFFSR_109 ( );
FILL FILL_47_DFFSR_109 ( );
FILL FILL_48_DFFSR_109 ( );
FILL FILL_49_DFFSR_109 ( );
FILL FILL_50_DFFSR_109 ( );
FILL FILL_0_DFFSR_96 ( );
FILL FILL_1_DFFSR_96 ( );
FILL FILL_2_DFFSR_96 ( );
FILL FILL_3_DFFSR_96 ( );
FILL FILL_4_DFFSR_96 ( );
FILL FILL_5_DFFSR_96 ( );
FILL FILL_6_DFFSR_96 ( );
FILL FILL_7_DFFSR_96 ( );
FILL FILL_8_DFFSR_96 ( );
FILL FILL_9_DFFSR_96 ( );
FILL FILL_10_DFFSR_96 ( );
FILL FILL_11_DFFSR_96 ( );
FILL FILL_12_DFFSR_96 ( );
FILL FILL_13_DFFSR_96 ( );
FILL FILL_14_DFFSR_96 ( );
FILL FILL_15_DFFSR_96 ( );
FILL FILL_16_DFFSR_96 ( );
FILL FILL_17_DFFSR_96 ( );
FILL FILL_18_DFFSR_96 ( );
FILL FILL_19_DFFSR_96 ( );
FILL FILL_20_DFFSR_96 ( );
FILL FILL_21_DFFSR_96 ( );
FILL FILL_22_DFFSR_96 ( );
FILL FILL_23_DFFSR_96 ( );
FILL FILL_24_DFFSR_96 ( );
FILL FILL_25_DFFSR_96 ( );
FILL FILL_26_DFFSR_96 ( );
FILL FILL_27_DFFSR_96 ( );
FILL FILL_28_DFFSR_96 ( );
FILL FILL_29_DFFSR_96 ( );
FILL FILL_30_DFFSR_96 ( );
FILL FILL_31_DFFSR_96 ( );
FILL FILL_32_DFFSR_96 ( );
FILL FILL_33_DFFSR_96 ( );
FILL FILL_34_DFFSR_96 ( );
FILL FILL_35_DFFSR_96 ( );
FILL FILL_36_DFFSR_96 ( );
FILL FILL_37_DFFSR_96 ( );
FILL FILL_38_DFFSR_96 ( );
FILL FILL_39_DFFSR_96 ( );
FILL FILL_40_DFFSR_96 ( );
FILL FILL_41_DFFSR_96 ( );
FILL FILL_42_DFFSR_96 ( );
FILL FILL_43_DFFSR_96 ( );
FILL FILL_44_DFFSR_96 ( );
FILL FILL_45_DFFSR_96 ( );
FILL FILL_46_DFFSR_96 ( );
FILL FILL_47_DFFSR_96 ( );
FILL FILL_48_DFFSR_96 ( );
FILL FILL_49_DFFSR_96 ( );
FILL FILL_50_DFFSR_96 ( );
FILL FILL_0_INVX1_185 ( );
FILL FILL_1_INVX1_185 ( );
FILL FILL_2_INVX1_185 ( );
FILL FILL_3_INVX1_185 ( );
FILL FILL_4_INVX1_185 ( );
FILL FILL_0_NAND3X1_231 ( );
FILL FILL_1_NAND3X1_231 ( );
FILL FILL_2_NAND3X1_231 ( );
FILL FILL_3_NAND3X1_231 ( );
FILL FILL_4_NAND3X1_231 ( );
FILL FILL_5_NAND3X1_231 ( );
FILL FILL_6_NAND3X1_231 ( );
FILL FILL_7_NAND3X1_231 ( );
FILL FILL_8_NAND3X1_231 ( );
FILL FILL_0_INVX1_173 ( );
FILL FILL_1_INVX1_173 ( );
FILL FILL_2_INVX1_173 ( );
FILL FILL_3_INVX1_173 ( );
FILL FILL_0_INVX1_178 ( );
FILL FILL_1_INVX1_178 ( );
FILL FILL_2_INVX1_178 ( );
FILL FILL_3_INVX1_178 ( );
FILL FILL_4_INVX1_178 ( );
FILL FILL_0_NAND3X1_236 ( );
FILL FILL_1_NAND3X1_236 ( );
FILL FILL_2_NAND3X1_236 ( );
FILL FILL_3_NAND3X1_236 ( );
FILL FILL_4_NAND3X1_236 ( );
FILL FILL_5_NAND3X1_236 ( );
FILL FILL_6_NAND3X1_236 ( );
FILL FILL_7_NAND3X1_236 ( );
FILL FILL_8_NAND3X1_236 ( );
FILL FILL_0_NAND3X1_232 ( );
FILL FILL_1_NAND3X1_232 ( );
FILL FILL_2_NAND3X1_232 ( );
FILL FILL_3_NAND3X1_232 ( );
FILL FILL_4_NAND3X1_232 ( );
FILL FILL_5_NAND3X1_232 ( );
FILL FILL_6_NAND3X1_232 ( );
FILL FILL_7_NAND3X1_232 ( );
FILL FILL_8_NAND3X1_232 ( );
FILL FILL_9_NAND3X1_232 ( );
FILL FILL_0_DFFSR_264 ( );
FILL FILL_1_DFFSR_264 ( );
FILL FILL_2_DFFSR_264 ( );
FILL FILL_3_DFFSR_264 ( );
FILL FILL_4_DFFSR_264 ( );
FILL FILL_5_DFFSR_264 ( );
FILL FILL_6_DFFSR_264 ( );
FILL FILL_7_DFFSR_264 ( );
FILL FILL_8_DFFSR_264 ( );
FILL FILL_9_DFFSR_264 ( );
FILL FILL_10_DFFSR_264 ( );
FILL FILL_11_DFFSR_264 ( );
FILL FILL_12_DFFSR_264 ( );
FILL FILL_13_DFFSR_264 ( );
FILL FILL_14_DFFSR_264 ( );
FILL FILL_15_DFFSR_264 ( );
FILL FILL_16_DFFSR_264 ( );
FILL FILL_17_DFFSR_264 ( );
FILL FILL_18_DFFSR_264 ( );
FILL FILL_19_DFFSR_264 ( );
FILL FILL_20_DFFSR_264 ( );
FILL FILL_21_DFFSR_264 ( );
FILL FILL_22_DFFSR_264 ( );
FILL FILL_23_DFFSR_264 ( );
FILL FILL_24_DFFSR_264 ( );
FILL FILL_25_DFFSR_264 ( );
FILL FILL_26_DFFSR_264 ( );
FILL FILL_27_DFFSR_264 ( );
FILL FILL_28_DFFSR_264 ( );
FILL FILL_29_DFFSR_264 ( );
FILL FILL_30_DFFSR_264 ( );
FILL FILL_31_DFFSR_264 ( );
FILL FILL_32_DFFSR_264 ( );
FILL FILL_33_DFFSR_264 ( );
FILL FILL_34_DFFSR_264 ( );
FILL FILL_35_DFFSR_264 ( );
FILL FILL_36_DFFSR_264 ( );
FILL FILL_37_DFFSR_264 ( );
FILL FILL_38_DFFSR_264 ( );
FILL FILL_39_DFFSR_264 ( );
FILL FILL_40_DFFSR_264 ( );
FILL FILL_41_DFFSR_264 ( );
FILL FILL_42_DFFSR_264 ( );
FILL FILL_43_DFFSR_264 ( );
FILL FILL_44_DFFSR_264 ( );
FILL FILL_45_DFFSR_264 ( );
FILL FILL_46_DFFSR_264 ( );
FILL FILL_47_DFFSR_264 ( );
FILL FILL_48_DFFSR_264 ( );
FILL FILL_49_DFFSR_264 ( );
FILL FILL_50_DFFSR_264 ( );
FILL FILL_51_DFFSR_264 ( );
FILL FILL_0_DFFSR_44 ( );
FILL FILL_1_DFFSR_44 ( );
FILL FILL_2_DFFSR_44 ( );
FILL FILL_3_DFFSR_44 ( );
FILL FILL_4_DFFSR_44 ( );
FILL FILL_5_DFFSR_44 ( );
FILL FILL_6_DFFSR_44 ( );
FILL FILL_7_DFFSR_44 ( );
FILL FILL_8_DFFSR_44 ( );
FILL FILL_9_DFFSR_44 ( );
FILL FILL_10_DFFSR_44 ( );
FILL FILL_11_DFFSR_44 ( );
FILL FILL_12_DFFSR_44 ( );
FILL FILL_13_DFFSR_44 ( );
FILL FILL_14_DFFSR_44 ( );
FILL FILL_15_DFFSR_44 ( );
FILL FILL_16_DFFSR_44 ( );
FILL FILL_17_DFFSR_44 ( );
FILL FILL_18_DFFSR_44 ( );
FILL FILL_19_DFFSR_44 ( );
FILL FILL_20_DFFSR_44 ( );
FILL FILL_21_DFFSR_44 ( );
FILL FILL_22_DFFSR_44 ( );
FILL FILL_23_DFFSR_44 ( );
FILL FILL_24_DFFSR_44 ( );
FILL FILL_25_DFFSR_44 ( );
FILL FILL_26_DFFSR_44 ( );
FILL FILL_27_DFFSR_44 ( );
FILL FILL_28_DFFSR_44 ( );
FILL FILL_29_DFFSR_44 ( );
FILL FILL_30_DFFSR_44 ( );
FILL FILL_31_DFFSR_44 ( );
FILL FILL_32_DFFSR_44 ( );
FILL FILL_33_DFFSR_44 ( );
FILL FILL_34_DFFSR_44 ( );
FILL FILL_35_DFFSR_44 ( );
FILL FILL_36_DFFSR_44 ( );
FILL FILL_37_DFFSR_44 ( );
FILL FILL_38_DFFSR_44 ( );
FILL FILL_39_DFFSR_44 ( );
FILL FILL_40_DFFSR_44 ( );
FILL FILL_41_DFFSR_44 ( );
FILL FILL_42_DFFSR_44 ( );
FILL FILL_43_DFFSR_44 ( );
FILL FILL_44_DFFSR_44 ( );
FILL FILL_45_DFFSR_44 ( );
FILL FILL_46_DFFSR_44 ( );
FILL FILL_47_DFFSR_44 ( );
FILL FILL_48_DFFSR_44 ( );
FILL FILL_49_DFFSR_44 ( );
FILL FILL_50_DFFSR_44 ( );
FILL FILL_0_DFFSR_63 ( );
FILL FILL_1_DFFSR_63 ( );
FILL FILL_2_DFFSR_63 ( );
FILL FILL_3_DFFSR_63 ( );
FILL FILL_4_DFFSR_63 ( );
FILL FILL_5_DFFSR_63 ( );
FILL FILL_6_DFFSR_63 ( );
FILL FILL_7_DFFSR_63 ( );
FILL FILL_8_DFFSR_63 ( );
FILL FILL_9_DFFSR_63 ( );
FILL FILL_10_DFFSR_63 ( );
FILL FILL_11_DFFSR_63 ( );
FILL FILL_12_DFFSR_63 ( );
FILL FILL_13_DFFSR_63 ( );
FILL FILL_14_DFFSR_63 ( );
FILL FILL_15_DFFSR_63 ( );
FILL FILL_16_DFFSR_63 ( );
FILL FILL_17_DFFSR_63 ( );
FILL FILL_18_DFFSR_63 ( );
FILL FILL_19_DFFSR_63 ( );
FILL FILL_20_DFFSR_63 ( );
FILL FILL_21_DFFSR_63 ( );
FILL FILL_22_DFFSR_63 ( );
FILL FILL_23_DFFSR_63 ( );
FILL FILL_24_DFFSR_63 ( );
FILL FILL_25_DFFSR_63 ( );
FILL FILL_26_DFFSR_63 ( );
FILL FILL_27_DFFSR_63 ( );
FILL FILL_28_DFFSR_63 ( );
FILL FILL_29_DFFSR_63 ( );
FILL FILL_30_DFFSR_63 ( );
FILL FILL_31_DFFSR_63 ( );
FILL FILL_32_DFFSR_63 ( );
FILL FILL_33_DFFSR_63 ( );
FILL FILL_34_DFFSR_63 ( );
FILL FILL_35_DFFSR_63 ( );
FILL FILL_36_DFFSR_63 ( );
FILL FILL_37_DFFSR_63 ( );
FILL FILL_38_DFFSR_63 ( );
FILL FILL_39_DFFSR_63 ( );
FILL FILL_40_DFFSR_63 ( );
FILL FILL_41_DFFSR_63 ( );
FILL FILL_42_DFFSR_63 ( );
FILL FILL_43_DFFSR_63 ( );
FILL FILL_44_DFFSR_63 ( );
FILL FILL_45_DFFSR_63 ( );
FILL FILL_46_DFFSR_63 ( );
FILL FILL_47_DFFSR_63 ( );
FILL FILL_48_DFFSR_63 ( );
FILL FILL_49_DFFSR_63 ( );
FILL FILL_50_DFFSR_63 ( );
FILL FILL_51_DFFSR_63 ( );
FILL FILL_0_INVX1_48 ( );
FILL FILL_1_INVX1_48 ( );
FILL FILL_2_INVX1_48 ( );
FILL FILL_3_INVX1_48 ( );
FILL FILL_4_INVX1_48 ( );
FILL FILL_0_OAI22X1_20 ( );
FILL FILL_1_OAI22X1_20 ( );
FILL FILL_2_OAI22X1_20 ( );
FILL FILL_3_OAI22X1_20 ( );
FILL FILL_4_OAI22X1_20 ( );
FILL FILL_5_OAI22X1_20 ( );
FILL FILL_6_OAI22X1_20 ( );
FILL FILL_7_OAI22X1_20 ( );
FILL FILL_8_OAI22X1_20 ( );
FILL FILL_9_OAI22X1_20 ( );
FILL FILL_10_OAI22X1_20 ( );
FILL FILL_11_OAI22X1_20 ( );
FILL FILL_0_OAI22X1_17 ( );
FILL FILL_1_OAI22X1_17 ( );
FILL FILL_2_OAI22X1_17 ( );
FILL FILL_3_OAI22X1_17 ( );
FILL FILL_4_OAI22X1_17 ( );
FILL FILL_5_OAI22X1_17 ( );
FILL FILL_6_OAI22X1_17 ( );
FILL FILL_7_OAI22X1_17 ( );
FILL FILL_8_OAI22X1_17 ( );
FILL FILL_9_OAI22X1_17 ( );
FILL FILL_10_OAI22X1_17 ( );
FILL FILL_11_OAI22X1_17 ( );
FILL FILL_0_INVX1_40 ( );
FILL FILL_1_INVX1_40 ( );
FILL FILL_2_INVX1_40 ( );
FILL FILL_3_INVX1_40 ( );
FILL FILL_4_INVX1_40 ( );
FILL FILL_0_INVX1_41 ( );
FILL FILL_1_INVX1_41 ( );
FILL FILL_2_INVX1_41 ( );
FILL FILL_3_INVX1_41 ( );
FILL FILL_0_OAI22X1_5 ( );
FILL FILL_1_OAI22X1_5 ( );
FILL FILL_2_OAI22X1_5 ( );
FILL FILL_3_OAI22X1_5 ( );
FILL FILL_4_OAI22X1_5 ( );
FILL FILL_5_OAI22X1_5 ( );
FILL FILL_6_OAI22X1_5 ( );
FILL FILL_7_OAI22X1_5 ( );
FILL FILL_8_OAI22X1_5 ( );
FILL FILL_9_OAI22X1_5 ( );
FILL FILL_10_OAI22X1_5 ( );
FILL FILL_11_OAI22X1_5 ( );
FILL FILL_0_INVX1_13 ( );
FILL FILL_1_INVX1_13 ( );
FILL FILL_2_INVX1_13 ( );
FILL FILL_3_INVX1_13 ( );
FILL FILL_4_INVX1_13 ( );
FILL FILL_0_DFFSR_102 ( );
FILL FILL_1_DFFSR_102 ( );
FILL FILL_2_DFFSR_102 ( );
FILL FILL_3_DFFSR_102 ( );
FILL FILL_4_DFFSR_102 ( );
FILL FILL_5_DFFSR_102 ( );
FILL FILL_6_DFFSR_102 ( );
FILL FILL_7_DFFSR_102 ( );
FILL FILL_8_DFFSR_102 ( );
FILL FILL_9_DFFSR_102 ( );
FILL FILL_10_DFFSR_102 ( );
FILL FILL_11_DFFSR_102 ( );
FILL FILL_12_DFFSR_102 ( );
FILL FILL_13_DFFSR_102 ( );
FILL FILL_14_DFFSR_102 ( );
FILL FILL_15_DFFSR_102 ( );
FILL FILL_16_DFFSR_102 ( );
FILL FILL_17_DFFSR_102 ( );
FILL FILL_18_DFFSR_102 ( );
FILL FILL_19_DFFSR_102 ( );
FILL FILL_20_DFFSR_102 ( );
FILL FILL_21_DFFSR_102 ( );
FILL FILL_22_DFFSR_102 ( );
FILL FILL_23_DFFSR_102 ( );
FILL FILL_24_DFFSR_102 ( );
FILL FILL_25_DFFSR_102 ( );
FILL FILL_26_DFFSR_102 ( );
FILL FILL_27_DFFSR_102 ( );
FILL FILL_28_DFFSR_102 ( );
FILL FILL_29_DFFSR_102 ( );
FILL FILL_30_DFFSR_102 ( );
FILL FILL_31_DFFSR_102 ( );
FILL FILL_32_DFFSR_102 ( );
FILL FILL_33_DFFSR_102 ( );
FILL FILL_34_DFFSR_102 ( );
FILL FILL_35_DFFSR_102 ( );
FILL FILL_36_DFFSR_102 ( );
FILL FILL_37_DFFSR_102 ( );
FILL FILL_38_DFFSR_102 ( );
FILL FILL_39_DFFSR_102 ( );
FILL FILL_40_DFFSR_102 ( );
FILL FILL_41_DFFSR_102 ( );
FILL FILL_42_DFFSR_102 ( );
FILL FILL_43_DFFSR_102 ( );
FILL FILL_44_DFFSR_102 ( );
FILL FILL_45_DFFSR_102 ( );
FILL FILL_46_DFFSR_102 ( );
FILL FILL_47_DFFSR_102 ( );
FILL FILL_48_DFFSR_102 ( );
FILL FILL_49_DFFSR_102 ( );
FILL FILL_50_DFFSR_102 ( );
FILL FILL_0_AOI22X1_2 ( );
FILL FILL_1_AOI22X1_2 ( );
FILL FILL_2_AOI22X1_2 ( );
FILL FILL_3_AOI22X1_2 ( );
FILL FILL_4_AOI22X1_2 ( );
FILL FILL_5_AOI22X1_2 ( );
FILL FILL_6_AOI22X1_2 ( );
FILL FILL_7_AOI22X1_2 ( );
FILL FILL_8_AOI22X1_2 ( );
FILL FILL_9_AOI22X1_2 ( );
FILL FILL_10_AOI22X1_2 ( );
FILL FILL_11_AOI22X1_2 ( );
FILL FILL_0_INVX1_55 ( );
FILL FILL_1_INVX1_55 ( );
FILL FILL_2_INVX1_55 ( );
FILL FILL_3_INVX1_55 ( );
FILL FILL_4_INVX1_55 ( );
FILL FILL_0_CLKBUF1_42 ( );
FILL FILL_1_CLKBUF1_42 ( );
FILL FILL_2_CLKBUF1_42 ( );
FILL FILL_3_CLKBUF1_42 ( );
FILL FILL_4_CLKBUF1_42 ( );
FILL FILL_5_CLKBUF1_42 ( );
FILL FILL_6_CLKBUF1_42 ( );
FILL FILL_7_CLKBUF1_42 ( );
FILL FILL_8_CLKBUF1_42 ( );
FILL FILL_9_CLKBUF1_42 ( );
FILL FILL_10_CLKBUF1_42 ( );
FILL FILL_11_CLKBUF1_42 ( );
FILL FILL_12_CLKBUF1_42 ( );
FILL FILL_13_CLKBUF1_42 ( );
FILL FILL_14_CLKBUF1_42 ( );
FILL FILL_15_CLKBUF1_42 ( );
FILL FILL_16_CLKBUF1_42 ( );
FILL FILL_17_CLKBUF1_42 ( );
FILL FILL_18_CLKBUF1_42 ( );
FILL FILL_19_CLKBUF1_42 ( );
FILL FILL_20_CLKBUF1_42 ( );
FILL FILL_0_CLKBUF1_24 ( );
FILL FILL_1_CLKBUF1_24 ( );
FILL FILL_2_CLKBUF1_24 ( );
FILL FILL_3_CLKBUF1_24 ( );
FILL FILL_4_CLKBUF1_24 ( );
FILL FILL_5_CLKBUF1_24 ( );
FILL FILL_6_CLKBUF1_24 ( );
FILL FILL_7_CLKBUF1_24 ( );
FILL FILL_8_CLKBUF1_24 ( );
FILL FILL_9_CLKBUF1_24 ( );
FILL FILL_10_CLKBUF1_24 ( );
FILL FILL_11_CLKBUF1_24 ( );
FILL FILL_12_CLKBUF1_24 ( );
FILL FILL_13_CLKBUF1_24 ( );
FILL FILL_14_CLKBUF1_24 ( );
FILL FILL_15_CLKBUF1_24 ( );
FILL FILL_16_CLKBUF1_24 ( );
FILL FILL_17_CLKBUF1_24 ( );
FILL FILL_18_CLKBUF1_24 ( );
FILL FILL_19_CLKBUF1_24 ( );
FILL FILL_20_CLKBUF1_24 ( );
FILL FILL_0_DFFSR_88 ( );
FILL FILL_1_DFFSR_88 ( );
FILL FILL_2_DFFSR_88 ( );
FILL FILL_3_DFFSR_88 ( );
FILL FILL_4_DFFSR_88 ( );
FILL FILL_5_DFFSR_88 ( );
FILL FILL_6_DFFSR_88 ( );
FILL FILL_7_DFFSR_88 ( );
FILL FILL_8_DFFSR_88 ( );
FILL FILL_9_DFFSR_88 ( );
FILL FILL_10_DFFSR_88 ( );
FILL FILL_11_DFFSR_88 ( );
FILL FILL_12_DFFSR_88 ( );
FILL FILL_13_DFFSR_88 ( );
FILL FILL_14_DFFSR_88 ( );
FILL FILL_15_DFFSR_88 ( );
FILL FILL_16_DFFSR_88 ( );
FILL FILL_17_DFFSR_88 ( );
FILL FILL_18_DFFSR_88 ( );
FILL FILL_19_DFFSR_88 ( );
FILL FILL_20_DFFSR_88 ( );
FILL FILL_21_DFFSR_88 ( );
FILL FILL_22_DFFSR_88 ( );
FILL FILL_23_DFFSR_88 ( );
FILL FILL_24_DFFSR_88 ( );
FILL FILL_25_DFFSR_88 ( );
FILL FILL_26_DFFSR_88 ( );
FILL FILL_27_DFFSR_88 ( );
FILL FILL_28_DFFSR_88 ( );
FILL FILL_29_DFFSR_88 ( );
FILL FILL_30_DFFSR_88 ( );
FILL FILL_31_DFFSR_88 ( );
FILL FILL_32_DFFSR_88 ( );
FILL FILL_33_DFFSR_88 ( );
FILL FILL_34_DFFSR_88 ( );
FILL FILL_35_DFFSR_88 ( );
FILL FILL_36_DFFSR_88 ( );
FILL FILL_37_DFFSR_88 ( );
FILL FILL_38_DFFSR_88 ( );
FILL FILL_39_DFFSR_88 ( );
FILL FILL_40_DFFSR_88 ( );
FILL FILL_41_DFFSR_88 ( );
FILL FILL_42_DFFSR_88 ( );
FILL FILL_43_DFFSR_88 ( );
FILL FILL_44_DFFSR_88 ( );
FILL FILL_45_DFFSR_88 ( );
FILL FILL_46_DFFSR_88 ( );
FILL FILL_47_DFFSR_88 ( );
FILL FILL_48_DFFSR_88 ( );
FILL FILL_49_DFFSR_88 ( );
FILL FILL_50_DFFSR_88 ( );
FILL FILL_0_CLKBUF1_23 ( );
FILL FILL_1_CLKBUF1_23 ( );
FILL FILL_2_CLKBUF1_23 ( );
FILL FILL_3_CLKBUF1_23 ( );
FILL FILL_4_CLKBUF1_23 ( );
FILL FILL_5_CLKBUF1_23 ( );
FILL FILL_6_CLKBUF1_23 ( );
FILL FILL_7_CLKBUF1_23 ( );
FILL FILL_8_CLKBUF1_23 ( );
FILL FILL_9_CLKBUF1_23 ( );
FILL FILL_10_CLKBUF1_23 ( );
FILL FILL_11_CLKBUF1_23 ( );
FILL FILL_12_CLKBUF1_23 ( );
FILL FILL_13_CLKBUF1_23 ( );
FILL FILL_14_CLKBUF1_23 ( );
FILL FILL_15_CLKBUF1_23 ( );
FILL FILL_16_CLKBUF1_23 ( );
FILL FILL_17_CLKBUF1_23 ( );
FILL FILL_18_CLKBUF1_23 ( );
FILL FILL_19_CLKBUF1_23 ( );
FILL FILL_0_DFFSR_226 ( );
FILL FILL_1_DFFSR_226 ( );
FILL FILL_2_DFFSR_226 ( );
FILL FILL_3_DFFSR_226 ( );
FILL FILL_4_DFFSR_226 ( );
FILL FILL_5_DFFSR_226 ( );
FILL FILL_6_DFFSR_226 ( );
FILL FILL_7_DFFSR_226 ( );
FILL FILL_8_DFFSR_226 ( );
FILL FILL_9_DFFSR_226 ( );
FILL FILL_10_DFFSR_226 ( );
FILL FILL_11_DFFSR_226 ( );
FILL FILL_12_DFFSR_226 ( );
FILL FILL_13_DFFSR_226 ( );
FILL FILL_14_DFFSR_226 ( );
FILL FILL_15_DFFSR_226 ( );
FILL FILL_16_DFFSR_226 ( );
FILL FILL_17_DFFSR_226 ( );
FILL FILL_18_DFFSR_226 ( );
FILL FILL_19_DFFSR_226 ( );
FILL FILL_20_DFFSR_226 ( );
FILL FILL_21_DFFSR_226 ( );
FILL FILL_22_DFFSR_226 ( );
FILL FILL_23_DFFSR_226 ( );
FILL FILL_24_DFFSR_226 ( );
FILL FILL_25_DFFSR_226 ( );
FILL FILL_26_DFFSR_226 ( );
FILL FILL_27_DFFSR_226 ( );
FILL FILL_28_DFFSR_226 ( );
FILL FILL_29_DFFSR_226 ( );
FILL FILL_30_DFFSR_226 ( );
FILL FILL_31_DFFSR_226 ( );
FILL FILL_32_DFFSR_226 ( );
FILL FILL_33_DFFSR_226 ( );
FILL FILL_34_DFFSR_226 ( );
FILL FILL_35_DFFSR_226 ( );
FILL FILL_36_DFFSR_226 ( );
FILL FILL_37_DFFSR_226 ( );
FILL FILL_38_DFFSR_226 ( );
FILL FILL_39_DFFSR_226 ( );
FILL FILL_40_DFFSR_226 ( );
FILL FILL_41_DFFSR_226 ( );
FILL FILL_42_DFFSR_226 ( );
FILL FILL_43_DFFSR_226 ( );
FILL FILL_44_DFFSR_226 ( );
FILL FILL_45_DFFSR_226 ( );
FILL FILL_46_DFFSR_226 ( );
FILL FILL_47_DFFSR_226 ( );
FILL FILL_48_DFFSR_226 ( );
FILL FILL_49_DFFSR_226 ( );
FILL FILL_50_DFFSR_226 ( );
FILL FILL_51_DFFSR_226 ( );
FILL FILL_0_AOI21X1_36 ( );
FILL FILL_1_AOI21X1_36 ( );
FILL FILL_2_AOI21X1_36 ( );
FILL FILL_3_AOI21X1_36 ( );
FILL FILL_4_AOI21X1_36 ( );
FILL FILL_5_AOI21X1_36 ( );
FILL FILL_6_AOI21X1_36 ( );
FILL FILL_7_AOI21X1_36 ( );
FILL FILL_8_AOI21X1_36 ( );
FILL FILL_9_AOI21X1_36 ( );
FILL FILL_0_NAND3X1_238 ( );
FILL FILL_1_NAND3X1_238 ( );
FILL FILL_2_NAND3X1_238 ( );
FILL FILL_3_NAND3X1_238 ( );
FILL FILL_4_NAND3X1_238 ( );
FILL FILL_5_NAND3X1_238 ( );
FILL FILL_6_NAND3X1_238 ( );
FILL FILL_7_NAND3X1_238 ( );
FILL FILL_8_NAND3X1_238 ( );
FILL FILL_0_NAND3X1_234 ( );
FILL FILL_1_NAND3X1_234 ( );
FILL FILL_2_NAND3X1_234 ( );
FILL FILL_3_NAND3X1_234 ( );
FILL FILL_4_NAND3X1_234 ( );
FILL FILL_5_NAND3X1_234 ( );
FILL FILL_6_NAND3X1_234 ( );
FILL FILL_7_NAND3X1_234 ( );
FILL FILL_8_NAND3X1_234 ( );
FILL FILL_0_DFFPOSX1_30 ( );
FILL FILL_1_DFFPOSX1_30 ( );
FILL FILL_2_DFFPOSX1_30 ( );
FILL FILL_3_DFFPOSX1_30 ( );
FILL FILL_4_DFFPOSX1_30 ( );
FILL FILL_5_DFFPOSX1_30 ( );
FILL FILL_6_DFFPOSX1_30 ( );
FILL FILL_7_DFFPOSX1_30 ( );
FILL FILL_8_DFFPOSX1_30 ( );
FILL FILL_9_DFFPOSX1_30 ( );
FILL FILL_10_DFFPOSX1_30 ( );
FILL FILL_11_DFFPOSX1_30 ( );
FILL FILL_12_DFFPOSX1_30 ( );
FILL FILL_13_DFFPOSX1_30 ( );
FILL FILL_14_DFFPOSX1_30 ( );
FILL FILL_15_DFFPOSX1_30 ( );
FILL FILL_16_DFFPOSX1_30 ( );
FILL FILL_17_DFFPOSX1_30 ( );
FILL FILL_18_DFFPOSX1_30 ( );
FILL FILL_19_DFFPOSX1_30 ( );
FILL FILL_20_DFFPOSX1_30 ( );
FILL FILL_21_DFFPOSX1_30 ( );
FILL FILL_22_DFFPOSX1_30 ( );
FILL FILL_23_DFFPOSX1_30 ( );
FILL FILL_24_DFFPOSX1_30 ( );
FILL FILL_25_DFFPOSX1_30 ( );
FILL FILL_26_DFFPOSX1_30 ( );
FILL FILL_27_DFFPOSX1_30 ( );
FILL FILL_0_INVX1_188 ( );
FILL FILL_1_INVX1_188 ( );
FILL FILL_2_INVX1_188 ( );
FILL FILL_3_INVX1_188 ( );
FILL FILL_4_INVX1_188 ( );
FILL FILL_0_OAI21X1_92 ( );
FILL FILL_1_OAI21X1_92 ( );
FILL FILL_2_OAI21X1_92 ( );
FILL FILL_3_OAI21X1_92 ( );
FILL FILL_4_OAI21X1_92 ( );
FILL FILL_5_OAI21X1_92 ( );
FILL FILL_6_OAI21X1_92 ( );
FILL FILL_7_OAI21X1_92 ( );
FILL FILL_8_OAI21X1_92 ( );
FILL FILL_0_NAND2X1_123 ( );
FILL FILL_1_NAND2X1_123 ( );
FILL FILL_2_NAND2X1_123 ( );
FILL FILL_3_NAND2X1_123 ( );
FILL FILL_4_NAND2X1_123 ( );
FILL FILL_5_NAND2X1_123 ( );
FILL FILL_6_NAND2X1_123 ( );
FILL FILL_0_DFFSR_36 ( );
FILL FILL_1_DFFSR_36 ( );
FILL FILL_2_DFFSR_36 ( );
FILL FILL_3_DFFSR_36 ( );
FILL FILL_4_DFFSR_36 ( );
FILL FILL_5_DFFSR_36 ( );
FILL FILL_6_DFFSR_36 ( );
FILL FILL_7_DFFSR_36 ( );
FILL FILL_8_DFFSR_36 ( );
FILL FILL_9_DFFSR_36 ( );
FILL FILL_10_DFFSR_36 ( );
FILL FILL_11_DFFSR_36 ( );
FILL FILL_12_DFFSR_36 ( );
FILL FILL_13_DFFSR_36 ( );
FILL FILL_14_DFFSR_36 ( );
FILL FILL_15_DFFSR_36 ( );
FILL FILL_16_DFFSR_36 ( );
FILL FILL_17_DFFSR_36 ( );
FILL FILL_18_DFFSR_36 ( );
FILL FILL_19_DFFSR_36 ( );
FILL FILL_20_DFFSR_36 ( );
FILL FILL_21_DFFSR_36 ( );
FILL FILL_22_DFFSR_36 ( );
FILL FILL_23_DFFSR_36 ( );
FILL FILL_24_DFFSR_36 ( );
FILL FILL_25_DFFSR_36 ( );
FILL FILL_26_DFFSR_36 ( );
FILL FILL_27_DFFSR_36 ( );
FILL FILL_28_DFFSR_36 ( );
FILL FILL_29_DFFSR_36 ( );
FILL FILL_30_DFFSR_36 ( );
FILL FILL_31_DFFSR_36 ( );
FILL FILL_32_DFFSR_36 ( );
FILL FILL_33_DFFSR_36 ( );
FILL FILL_34_DFFSR_36 ( );
FILL FILL_35_DFFSR_36 ( );
FILL FILL_36_DFFSR_36 ( );
FILL FILL_37_DFFSR_36 ( );
FILL FILL_38_DFFSR_36 ( );
FILL FILL_39_DFFSR_36 ( );
FILL FILL_40_DFFSR_36 ( );
FILL FILL_41_DFFSR_36 ( );
FILL FILL_42_DFFSR_36 ( );
FILL FILL_43_DFFSR_36 ( );
FILL FILL_44_DFFSR_36 ( );
FILL FILL_45_DFFSR_36 ( );
FILL FILL_46_DFFSR_36 ( );
FILL FILL_47_DFFSR_36 ( );
FILL FILL_48_DFFSR_36 ( );
FILL FILL_49_DFFSR_36 ( );
FILL FILL_50_DFFSR_36 ( );
FILL FILL_51_DFFSR_36 ( );
FILL FILL_0_DFFSR_47 ( );
FILL FILL_1_DFFSR_47 ( );
FILL FILL_2_DFFSR_47 ( );
FILL FILL_3_DFFSR_47 ( );
FILL FILL_4_DFFSR_47 ( );
FILL FILL_5_DFFSR_47 ( );
FILL FILL_6_DFFSR_47 ( );
FILL FILL_7_DFFSR_47 ( );
FILL FILL_8_DFFSR_47 ( );
FILL FILL_9_DFFSR_47 ( );
FILL FILL_10_DFFSR_47 ( );
FILL FILL_11_DFFSR_47 ( );
FILL FILL_12_DFFSR_47 ( );
FILL FILL_13_DFFSR_47 ( );
FILL FILL_14_DFFSR_47 ( );
FILL FILL_15_DFFSR_47 ( );
FILL FILL_16_DFFSR_47 ( );
FILL FILL_17_DFFSR_47 ( );
FILL FILL_18_DFFSR_47 ( );
FILL FILL_19_DFFSR_47 ( );
FILL FILL_20_DFFSR_47 ( );
FILL FILL_21_DFFSR_47 ( );
FILL FILL_22_DFFSR_47 ( );
FILL FILL_23_DFFSR_47 ( );
FILL FILL_24_DFFSR_47 ( );
FILL FILL_25_DFFSR_47 ( );
FILL FILL_26_DFFSR_47 ( );
FILL FILL_27_DFFSR_47 ( );
FILL FILL_28_DFFSR_47 ( );
FILL FILL_29_DFFSR_47 ( );
FILL FILL_30_DFFSR_47 ( );
FILL FILL_31_DFFSR_47 ( );
FILL FILL_32_DFFSR_47 ( );
FILL FILL_33_DFFSR_47 ( );
FILL FILL_34_DFFSR_47 ( );
FILL FILL_35_DFFSR_47 ( );
FILL FILL_36_DFFSR_47 ( );
FILL FILL_37_DFFSR_47 ( );
FILL FILL_38_DFFSR_47 ( );
FILL FILL_39_DFFSR_47 ( );
FILL FILL_40_DFFSR_47 ( );
FILL FILL_41_DFFSR_47 ( );
FILL FILL_42_DFFSR_47 ( );
FILL FILL_43_DFFSR_47 ( );
FILL FILL_44_DFFSR_47 ( );
FILL FILL_45_DFFSR_47 ( );
FILL FILL_46_DFFSR_47 ( );
FILL FILL_47_DFFSR_47 ( );
FILL FILL_48_DFFSR_47 ( );
FILL FILL_49_DFFSR_47 ( );
FILL FILL_50_DFFSR_47 ( );
FILL FILL_0_INVX1_47 ( );
FILL FILL_1_INVX1_47 ( );
FILL FILL_2_INVX1_47 ( );
FILL FILL_3_INVX1_47 ( );
FILL FILL_0_DFFSR_94 ( );
FILL FILL_1_DFFSR_94 ( );
FILL FILL_2_DFFSR_94 ( );
FILL FILL_3_DFFSR_94 ( );
FILL FILL_4_DFFSR_94 ( );
FILL FILL_5_DFFSR_94 ( );
FILL FILL_6_DFFSR_94 ( );
FILL FILL_7_DFFSR_94 ( );
FILL FILL_8_DFFSR_94 ( );
FILL FILL_9_DFFSR_94 ( );
FILL FILL_10_DFFSR_94 ( );
FILL FILL_11_DFFSR_94 ( );
FILL FILL_12_DFFSR_94 ( );
FILL FILL_13_DFFSR_94 ( );
FILL FILL_14_DFFSR_94 ( );
FILL FILL_15_DFFSR_94 ( );
FILL FILL_16_DFFSR_94 ( );
FILL FILL_17_DFFSR_94 ( );
FILL FILL_18_DFFSR_94 ( );
FILL FILL_19_DFFSR_94 ( );
FILL FILL_20_DFFSR_94 ( );
FILL FILL_21_DFFSR_94 ( );
FILL FILL_22_DFFSR_94 ( );
FILL FILL_23_DFFSR_94 ( );
FILL FILL_24_DFFSR_94 ( );
FILL FILL_25_DFFSR_94 ( );
FILL FILL_26_DFFSR_94 ( );
FILL FILL_27_DFFSR_94 ( );
FILL FILL_28_DFFSR_94 ( );
FILL FILL_29_DFFSR_94 ( );
FILL FILL_30_DFFSR_94 ( );
FILL FILL_31_DFFSR_94 ( );
FILL FILL_32_DFFSR_94 ( );
FILL FILL_33_DFFSR_94 ( );
FILL FILL_34_DFFSR_94 ( );
FILL FILL_35_DFFSR_94 ( );
FILL FILL_36_DFFSR_94 ( );
FILL FILL_37_DFFSR_94 ( );
FILL FILL_38_DFFSR_94 ( );
FILL FILL_39_DFFSR_94 ( );
FILL FILL_40_DFFSR_94 ( );
FILL FILL_41_DFFSR_94 ( );
FILL FILL_42_DFFSR_94 ( );
FILL FILL_43_DFFSR_94 ( );
FILL FILL_44_DFFSR_94 ( );
FILL FILL_45_DFFSR_94 ( );
FILL FILL_46_DFFSR_94 ( );
FILL FILL_47_DFFSR_94 ( );
FILL FILL_48_DFFSR_94 ( );
FILL FILL_49_DFFSR_94 ( );
FILL FILL_50_DFFSR_94 ( );
FILL FILL_0_DFFSR_82 ( );
FILL FILL_1_DFFSR_82 ( );
FILL FILL_2_DFFSR_82 ( );
FILL FILL_3_DFFSR_82 ( );
FILL FILL_4_DFFSR_82 ( );
FILL FILL_5_DFFSR_82 ( );
FILL FILL_6_DFFSR_82 ( );
FILL FILL_7_DFFSR_82 ( );
FILL FILL_8_DFFSR_82 ( );
FILL FILL_9_DFFSR_82 ( );
FILL FILL_10_DFFSR_82 ( );
FILL FILL_11_DFFSR_82 ( );
FILL FILL_12_DFFSR_82 ( );
FILL FILL_13_DFFSR_82 ( );
FILL FILL_14_DFFSR_82 ( );
FILL FILL_15_DFFSR_82 ( );
FILL FILL_16_DFFSR_82 ( );
FILL FILL_17_DFFSR_82 ( );
FILL FILL_18_DFFSR_82 ( );
FILL FILL_19_DFFSR_82 ( );
FILL FILL_20_DFFSR_82 ( );
FILL FILL_21_DFFSR_82 ( );
FILL FILL_22_DFFSR_82 ( );
FILL FILL_23_DFFSR_82 ( );
FILL FILL_24_DFFSR_82 ( );
FILL FILL_25_DFFSR_82 ( );
FILL FILL_26_DFFSR_82 ( );
FILL FILL_27_DFFSR_82 ( );
FILL FILL_28_DFFSR_82 ( );
FILL FILL_29_DFFSR_82 ( );
FILL FILL_30_DFFSR_82 ( );
FILL FILL_31_DFFSR_82 ( );
FILL FILL_32_DFFSR_82 ( );
FILL FILL_33_DFFSR_82 ( );
FILL FILL_34_DFFSR_82 ( );
FILL FILL_35_DFFSR_82 ( );
FILL FILL_36_DFFSR_82 ( );
FILL FILL_37_DFFSR_82 ( );
FILL FILL_38_DFFSR_82 ( );
FILL FILL_39_DFFSR_82 ( );
FILL FILL_40_DFFSR_82 ( );
FILL FILL_41_DFFSR_82 ( );
FILL FILL_42_DFFSR_82 ( );
FILL FILL_43_DFFSR_82 ( );
FILL FILL_44_DFFSR_82 ( );
FILL FILL_45_DFFSR_82 ( );
FILL FILL_46_DFFSR_82 ( );
FILL FILL_47_DFFSR_82 ( );
FILL FILL_48_DFFSR_82 ( );
FILL FILL_49_DFFSR_82 ( );
FILL FILL_50_DFFSR_82 ( );
FILL FILL_0_DFFSR_98 ( );
FILL FILL_1_DFFSR_98 ( );
FILL FILL_2_DFFSR_98 ( );
FILL FILL_3_DFFSR_98 ( );
FILL FILL_4_DFFSR_98 ( );
FILL FILL_5_DFFSR_98 ( );
FILL FILL_6_DFFSR_98 ( );
FILL FILL_7_DFFSR_98 ( );
FILL FILL_8_DFFSR_98 ( );
FILL FILL_9_DFFSR_98 ( );
FILL FILL_10_DFFSR_98 ( );
FILL FILL_11_DFFSR_98 ( );
FILL FILL_12_DFFSR_98 ( );
FILL FILL_13_DFFSR_98 ( );
FILL FILL_14_DFFSR_98 ( );
FILL FILL_15_DFFSR_98 ( );
FILL FILL_16_DFFSR_98 ( );
FILL FILL_17_DFFSR_98 ( );
FILL FILL_18_DFFSR_98 ( );
FILL FILL_19_DFFSR_98 ( );
FILL FILL_20_DFFSR_98 ( );
FILL FILL_21_DFFSR_98 ( );
FILL FILL_22_DFFSR_98 ( );
FILL FILL_23_DFFSR_98 ( );
FILL FILL_24_DFFSR_98 ( );
FILL FILL_25_DFFSR_98 ( );
FILL FILL_26_DFFSR_98 ( );
FILL FILL_27_DFFSR_98 ( );
FILL FILL_28_DFFSR_98 ( );
FILL FILL_29_DFFSR_98 ( );
FILL FILL_30_DFFSR_98 ( );
FILL FILL_31_DFFSR_98 ( );
FILL FILL_32_DFFSR_98 ( );
FILL FILL_33_DFFSR_98 ( );
FILL FILL_34_DFFSR_98 ( );
FILL FILL_35_DFFSR_98 ( );
FILL FILL_36_DFFSR_98 ( );
FILL FILL_37_DFFSR_98 ( );
FILL FILL_38_DFFSR_98 ( );
FILL FILL_39_DFFSR_98 ( );
FILL FILL_40_DFFSR_98 ( );
FILL FILL_41_DFFSR_98 ( );
FILL FILL_42_DFFSR_98 ( );
FILL FILL_43_DFFSR_98 ( );
FILL FILL_44_DFFSR_98 ( );
FILL FILL_45_DFFSR_98 ( );
FILL FILL_46_DFFSR_98 ( );
FILL FILL_47_DFFSR_98 ( );
FILL FILL_48_DFFSR_98 ( );
FILL FILL_49_DFFSR_98 ( );
FILL FILL_50_DFFSR_98 ( );
FILL FILL_51_DFFSR_98 ( );
FILL FILL_0_INVX1_37 ( );
FILL FILL_1_INVX1_37 ( );
FILL FILL_2_INVX1_37 ( );
FILL FILL_3_INVX1_37 ( );
FILL FILL_4_INVX1_37 ( );
FILL FILL_0_DFFSR_117 ( );
FILL FILL_1_DFFSR_117 ( );
FILL FILL_2_DFFSR_117 ( );
FILL FILL_3_DFFSR_117 ( );
FILL FILL_4_DFFSR_117 ( );
FILL FILL_5_DFFSR_117 ( );
FILL FILL_6_DFFSR_117 ( );
FILL FILL_7_DFFSR_117 ( );
FILL FILL_8_DFFSR_117 ( );
FILL FILL_9_DFFSR_117 ( );
FILL FILL_10_DFFSR_117 ( );
FILL FILL_11_DFFSR_117 ( );
FILL FILL_12_DFFSR_117 ( );
FILL FILL_13_DFFSR_117 ( );
FILL FILL_14_DFFSR_117 ( );
FILL FILL_15_DFFSR_117 ( );
FILL FILL_16_DFFSR_117 ( );
FILL FILL_17_DFFSR_117 ( );
FILL FILL_18_DFFSR_117 ( );
FILL FILL_19_DFFSR_117 ( );
FILL FILL_20_DFFSR_117 ( );
FILL FILL_21_DFFSR_117 ( );
FILL FILL_22_DFFSR_117 ( );
FILL FILL_23_DFFSR_117 ( );
FILL FILL_24_DFFSR_117 ( );
FILL FILL_25_DFFSR_117 ( );
FILL FILL_26_DFFSR_117 ( );
FILL FILL_27_DFFSR_117 ( );
FILL FILL_28_DFFSR_117 ( );
FILL FILL_29_DFFSR_117 ( );
FILL FILL_30_DFFSR_117 ( );
FILL FILL_31_DFFSR_117 ( );
FILL FILL_32_DFFSR_117 ( );
FILL FILL_33_DFFSR_117 ( );
FILL FILL_34_DFFSR_117 ( );
FILL FILL_35_DFFSR_117 ( );
FILL FILL_36_DFFSR_117 ( );
FILL FILL_37_DFFSR_117 ( );
FILL FILL_38_DFFSR_117 ( );
FILL FILL_39_DFFSR_117 ( );
FILL FILL_40_DFFSR_117 ( );
FILL FILL_41_DFFSR_117 ( );
FILL FILL_42_DFFSR_117 ( );
FILL FILL_43_DFFSR_117 ( );
FILL FILL_44_DFFSR_117 ( );
FILL FILL_45_DFFSR_117 ( );
FILL FILL_46_DFFSR_117 ( );
FILL FILL_47_DFFSR_117 ( );
FILL FILL_48_DFFSR_117 ( );
FILL FILL_49_DFFSR_117 ( );
FILL FILL_50_DFFSR_117 ( );
FILL FILL_51_DFFSR_117 ( );
FILL FILL_0_DFFSR_261 ( );
FILL FILL_1_DFFSR_261 ( );
FILL FILL_2_DFFSR_261 ( );
FILL FILL_3_DFFSR_261 ( );
FILL FILL_4_DFFSR_261 ( );
FILL FILL_5_DFFSR_261 ( );
FILL FILL_6_DFFSR_261 ( );
FILL FILL_7_DFFSR_261 ( );
FILL FILL_8_DFFSR_261 ( );
FILL FILL_9_DFFSR_261 ( );
FILL FILL_10_DFFSR_261 ( );
FILL FILL_11_DFFSR_261 ( );
FILL FILL_12_DFFSR_261 ( );
FILL FILL_13_DFFSR_261 ( );
FILL FILL_14_DFFSR_261 ( );
FILL FILL_15_DFFSR_261 ( );
FILL FILL_16_DFFSR_261 ( );
FILL FILL_17_DFFSR_261 ( );
FILL FILL_18_DFFSR_261 ( );
FILL FILL_19_DFFSR_261 ( );
FILL FILL_20_DFFSR_261 ( );
FILL FILL_21_DFFSR_261 ( );
FILL FILL_22_DFFSR_261 ( );
FILL FILL_23_DFFSR_261 ( );
FILL FILL_24_DFFSR_261 ( );
FILL FILL_25_DFFSR_261 ( );
FILL FILL_26_DFFSR_261 ( );
FILL FILL_27_DFFSR_261 ( );
FILL FILL_28_DFFSR_261 ( );
FILL FILL_29_DFFSR_261 ( );
FILL FILL_30_DFFSR_261 ( );
FILL FILL_31_DFFSR_261 ( );
FILL FILL_32_DFFSR_261 ( );
FILL FILL_33_DFFSR_261 ( );
FILL FILL_34_DFFSR_261 ( );
FILL FILL_35_DFFSR_261 ( );
FILL FILL_36_DFFSR_261 ( );
FILL FILL_37_DFFSR_261 ( );
FILL FILL_38_DFFSR_261 ( );
FILL FILL_39_DFFSR_261 ( );
FILL FILL_40_DFFSR_261 ( );
FILL FILL_41_DFFSR_261 ( );
FILL FILL_42_DFFSR_261 ( );
FILL FILL_43_DFFSR_261 ( );
FILL FILL_44_DFFSR_261 ( );
FILL FILL_45_DFFSR_261 ( );
FILL FILL_46_DFFSR_261 ( );
FILL FILL_47_DFFSR_261 ( );
FILL FILL_48_DFFSR_261 ( );
FILL FILL_49_DFFSR_261 ( );
FILL FILL_50_DFFSR_261 ( );
FILL FILL_51_DFFSR_261 ( );
FILL FILL_0_NAND3X1_125 ( );
FILL FILL_1_NAND3X1_125 ( );
FILL FILL_2_NAND3X1_125 ( );
FILL FILL_3_NAND3X1_125 ( );
FILL FILL_4_NAND3X1_125 ( );
FILL FILL_5_NAND3X1_125 ( );
FILL FILL_6_NAND3X1_125 ( );
FILL FILL_7_NAND3X1_125 ( );
FILL FILL_8_NAND3X1_125 ( );
FILL FILL_0_BUFX2_86 ( );
FILL FILL_1_BUFX2_86 ( );
FILL FILL_2_BUFX2_86 ( );
FILL FILL_3_BUFX2_86 ( );
FILL FILL_4_BUFX2_86 ( );
FILL FILL_5_BUFX2_86 ( );
FILL FILL_6_BUFX2_86 ( );
FILL FILL_0_INVX1_113 ( );
FILL FILL_1_INVX1_113 ( );
FILL FILL_2_INVX1_113 ( );
FILL FILL_3_INVX1_113 ( );
FILL FILL_4_INVX1_113 ( );
FILL FILL_0_INVX1_96 ( );
FILL FILL_1_INVX1_96 ( );
FILL FILL_2_INVX1_96 ( );
FILL FILL_3_INVX1_96 ( );
FILL FILL_4_INVX1_96 ( );
FILL FILL_0_INVX1_114 ( );
FILL FILL_1_INVX1_114 ( );
FILL FILL_2_INVX1_114 ( );
FILL FILL_3_INVX1_114 ( );
FILL FILL_4_INVX1_114 ( );
FILL FILL_0_NAND2X1_117 ( );
FILL FILL_1_NAND2X1_117 ( );
FILL FILL_2_NAND2X1_117 ( );
FILL FILL_3_NAND2X1_117 ( );
FILL FILL_4_NAND2X1_117 ( );
FILL FILL_5_NAND2X1_117 ( );
FILL FILL_6_NAND2X1_117 ( );
FILL FILL_0_OAI21X1_86 ( );
FILL FILL_1_OAI21X1_86 ( );
FILL FILL_2_OAI21X1_86 ( );
FILL FILL_3_OAI21X1_86 ( );
FILL FILL_4_OAI21X1_86 ( );
FILL FILL_5_OAI21X1_86 ( );
FILL FILL_6_OAI21X1_86 ( );
FILL FILL_7_OAI21X1_86 ( );
FILL FILL_8_OAI21X1_86 ( );
FILL FILL_0_INVX1_182 ( );
FILL FILL_1_INVX1_182 ( );
FILL FILL_2_INVX1_182 ( );
FILL FILL_3_INVX1_182 ( );
FILL FILL_4_INVX1_182 ( );
FILL FILL_0_DFFSR_260 ( );
FILL FILL_1_DFFSR_260 ( );
FILL FILL_2_DFFSR_260 ( );
FILL FILL_3_DFFSR_260 ( );
FILL FILL_4_DFFSR_260 ( );
FILL FILL_5_DFFSR_260 ( );
FILL FILL_6_DFFSR_260 ( );
FILL FILL_7_DFFSR_260 ( );
FILL FILL_8_DFFSR_260 ( );
FILL FILL_9_DFFSR_260 ( );
FILL FILL_10_DFFSR_260 ( );
FILL FILL_11_DFFSR_260 ( );
FILL FILL_12_DFFSR_260 ( );
FILL FILL_13_DFFSR_260 ( );
FILL FILL_14_DFFSR_260 ( );
FILL FILL_15_DFFSR_260 ( );
FILL FILL_16_DFFSR_260 ( );
FILL FILL_17_DFFSR_260 ( );
FILL FILL_18_DFFSR_260 ( );
FILL FILL_19_DFFSR_260 ( );
FILL FILL_20_DFFSR_260 ( );
FILL FILL_21_DFFSR_260 ( );
FILL FILL_22_DFFSR_260 ( );
FILL FILL_23_DFFSR_260 ( );
FILL FILL_24_DFFSR_260 ( );
FILL FILL_25_DFFSR_260 ( );
FILL FILL_26_DFFSR_260 ( );
FILL FILL_27_DFFSR_260 ( );
FILL FILL_28_DFFSR_260 ( );
FILL FILL_29_DFFSR_260 ( );
FILL FILL_30_DFFSR_260 ( );
FILL FILL_31_DFFSR_260 ( );
FILL FILL_32_DFFSR_260 ( );
FILL FILL_33_DFFSR_260 ( );
FILL FILL_34_DFFSR_260 ( );
FILL FILL_35_DFFSR_260 ( );
FILL FILL_36_DFFSR_260 ( );
FILL FILL_37_DFFSR_260 ( );
FILL FILL_38_DFFSR_260 ( );
FILL FILL_39_DFFSR_260 ( );
FILL FILL_40_DFFSR_260 ( );
FILL FILL_41_DFFSR_260 ( );
FILL FILL_42_DFFSR_260 ( );
FILL FILL_43_DFFSR_260 ( );
FILL FILL_44_DFFSR_260 ( );
FILL FILL_45_DFFSR_260 ( );
FILL FILL_46_DFFSR_260 ( );
FILL FILL_47_DFFSR_260 ( );
FILL FILL_48_DFFSR_260 ( );
FILL FILL_49_DFFSR_260 ( );
FILL FILL_50_DFFSR_260 ( );
FILL FILL_0_BUFX2_77 ( );
FILL FILL_1_BUFX2_77 ( );
FILL FILL_2_BUFX2_77 ( );
FILL FILL_3_BUFX2_77 ( );
FILL FILL_4_BUFX2_77 ( );
FILL FILL_5_BUFX2_77 ( );
FILL FILL_6_BUFX2_77 ( );
FILL FILL_0_DFFSR_50 ( );
FILL FILL_1_DFFSR_50 ( );
FILL FILL_2_DFFSR_50 ( );
FILL FILL_3_DFFSR_50 ( );
FILL FILL_4_DFFSR_50 ( );
FILL FILL_5_DFFSR_50 ( );
FILL FILL_6_DFFSR_50 ( );
FILL FILL_7_DFFSR_50 ( );
FILL FILL_8_DFFSR_50 ( );
FILL FILL_9_DFFSR_50 ( );
FILL FILL_10_DFFSR_50 ( );
FILL FILL_11_DFFSR_50 ( );
FILL FILL_12_DFFSR_50 ( );
FILL FILL_13_DFFSR_50 ( );
FILL FILL_14_DFFSR_50 ( );
FILL FILL_15_DFFSR_50 ( );
FILL FILL_16_DFFSR_50 ( );
FILL FILL_17_DFFSR_50 ( );
FILL FILL_18_DFFSR_50 ( );
FILL FILL_19_DFFSR_50 ( );
FILL FILL_20_DFFSR_50 ( );
FILL FILL_21_DFFSR_50 ( );
FILL FILL_22_DFFSR_50 ( );
FILL FILL_23_DFFSR_50 ( );
FILL FILL_24_DFFSR_50 ( );
FILL FILL_25_DFFSR_50 ( );
FILL FILL_26_DFFSR_50 ( );
FILL FILL_27_DFFSR_50 ( );
FILL FILL_28_DFFSR_50 ( );
FILL FILL_29_DFFSR_50 ( );
FILL FILL_30_DFFSR_50 ( );
FILL FILL_31_DFFSR_50 ( );
FILL FILL_32_DFFSR_50 ( );
FILL FILL_33_DFFSR_50 ( );
FILL FILL_34_DFFSR_50 ( );
FILL FILL_35_DFFSR_50 ( );
FILL FILL_36_DFFSR_50 ( );
FILL FILL_37_DFFSR_50 ( );
FILL FILL_38_DFFSR_50 ( );
FILL FILL_39_DFFSR_50 ( );
FILL FILL_40_DFFSR_50 ( );
FILL FILL_41_DFFSR_50 ( );
FILL FILL_42_DFFSR_50 ( );
FILL FILL_43_DFFSR_50 ( );
FILL FILL_44_DFFSR_50 ( );
FILL FILL_45_DFFSR_50 ( );
FILL FILL_46_DFFSR_50 ( );
FILL FILL_47_DFFSR_50 ( );
FILL FILL_48_DFFSR_50 ( );
FILL FILL_49_DFFSR_50 ( );
FILL FILL_50_DFFSR_50 ( );
FILL FILL_0_BUFX2_50 ( );
FILL FILL_1_BUFX2_50 ( );
FILL FILL_2_BUFX2_50 ( );
FILL FILL_3_BUFX2_50 ( );
FILL FILL_4_BUFX2_50 ( );
FILL FILL_5_BUFX2_50 ( );
FILL FILL_6_BUFX2_50 ( );
FILL FILL_0_BUFX2_45 ( );
FILL FILL_1_BUFX2_45 ( );
FILL FILL_2_BUFX2_45 ( );
FILL FILL_3_BUFX2_45 ( );
FILL FILL_4_BUFX2_45 ( );
FILL FILL_5_BUFX2_45 ( );
FILL FILL_6_BUFX2_45 ( );
FILL FILL_0_INVX1_10 ( );
FILL FILL_1_INVX1_10 ( );
FILL FILL_2_INVX1_10 ( );
FILL FILL_3_INVX1_10 ( );
FILL FILL_0_DFFSR_87 ( );
FILL FILL_1_DFFSR_87 ( );
FILL FILL_2_DFFSR_87 ( );
FILL FILL_3_DFFSR_87 ( );
FILL FILL_4_DFFSR_87 ( );
FILL FILL_5_DFFSR_87 ( );
FILL FILL_6_DFFSR_87 ( );
FILL FILL_7_DFFSR_87 ( );
FILL FILL_8_DFFSR_87 ( );
FILL FILL_9_DFFSR_87 ( );
FILL FILL_10_DFFSR_87 ( );
FILL FILL_11_DFFSR_87 ( );
FILL FILL_12_DFFSR_87 ( );
FILL FILL_13_DFFSR_87 ( );
FILL FILL_14_DFFSR_87 ( );
FILL FILL_15_DFFSR_87 ( );
FILL FILL_16_DFFSR_87 ( );
FILL FILL_17_DFFSR_87 ( );
FILL FILL_18_DFFSR_87 ( );
FILL FILL_19_DFFSR_87 ( );
FILL FILL_20_DFFSR_87 ( );
FILL FILL_21_DFFSR_87 ( );
FILL FILL_22_DFFSR_87 ( );
FILL FILL_23_DFFSR_87 ( );
FILL FILL_24_DFFSR_87 ( );
FILL FILL_25_DFFSR_87 ( );
FILL FILL_26_DFFSR_87 ( );
FILL FILL_27_DFFSR_87 ( );
FILL FILL_28_DFFSR_87 ( );
FILL FILL_29_DFFSR_87 ( );
FILL FILL_30_DFFSR_87 ( );
FILL FILL_31_DFFSR_87 ( );
FILL FILL_32_DFFSR_87 ( );
FILL FILL_33_DFFSR_87 ( );
FILL FILL_34_DFFSR_87 ( );
FILL FILL_35_DFFSR_87 ( );
FILL FILL_36_DFFSR_87 ( );
FILL FILL_37_DFFSR_87 ( );
FILL FILL_38_DFFSR_87 ( );
FILL FILL_39_DFFSR_87 ( );
FILL FILL_40_DFFSR_87 ( );
FILL FILL_41_DFFSR_87 ( );
FILL FILL_42_DFFSR_87 ( );
FILL FILL_43_DFFSR_87 ( );
FILL FILL_44_DFFSR_87 ( );
FILL FILL_45_DFFSR_87 ( );
FILL FILL_46_DFFSR_87 ( );
FILL FILL_47_DFFSR_87 ( );
FILL FILL_48_DFFSR_87 ( );
FILL FILL_49_DFFSR_87 ( );
FILL FILL_50_DFFSR_87 ( );
FILL FILL_0_DFFSR_66 ( );
FILL FILL_1_DFFSR_66 ( );
FILL FILL_2_DFFSR_66 ( );
FILL FILL_3_DFFSR_66 ( );
FILL FILL_4_DFFSR_66 ( );
FILL FILL_5_DFFSR_66 ( );
FILL FILL_6_DFFSR_66 ( );
FILL FILL_7_DFFSR_66 ( );
FILL FILL_8_DFFSR_66 ( );
FILL FILL_9_DFFSR_66 ( );
FILL FILL_10_DFFSR_66 ( );
FILL FILL_11_DFFSR_66 ( );
FILL FILL_12_DFFSR_66 ( );
FILL FILL_13_DFFSR_66 ( );
FILL FILL_14_DFFSR_66 ( );
FILL FILL_15_DFFSR_66 ( );
FILL FILL_16_DFFSR_66 ( );
FILL FILL_17_DFFSR_66 ( );
FILL FILL_18_DFFSR_66 ( );
FILL FILL_19_DFFSR_66 ( );
FILL FILL_20_DFFSR_66 ( );
FILL FILL_21_DFFSR_66 ( );
FILL FILL_22_DFFSR_66 ( );
FILL FILL_23_DFFSR_66 ( );
FILL FILL_24_DFFSR_66 ( );
FILL FILL_25_DFFSR_66 ( );
FILL FILL_26_DFFSR_66 ( );
FILL FILL_27_DFFSR_66 ( );
FILL FILL_28_DFFSR_66 ( );
FILL FILL_29_DFFSR_66 ( );
FILL FILL_30_DFFSR_66 ( );
FILL FILL_31_DFFSR_66 ( );
FILL FILL_32_DFFSR_66 ( );
FILL FILL_33_DFFSR_66 ( );
FILL FILL_34_DFFSR_66 ( );
FILL FILL_35_DFFSR_66 ( );
FILL FILL_36_DFFSR_66 ( );
FILL FILL_37_DFFSR_66 ( );
FILL FILL_38_DFFSR_66 ( );
FILL FILL_39_DFFSR_66 ( );
FILL FILL_40_DFFSR_66 ( );
FILL FILL_41_DFFSR_66 ( );
FILL FILL_42_DFFSR_66 ( );
FILL FILL_43_DFFSR_66 ( );
FILL FILL_44_DFFSR_66 ( );
FILL FILL_45_DFFSR_66 ( );
FILL FILL_46_DFFSR_66 ( );
FILL FILL_47_DFFSR_66 ( );
FILL FILL_48_DFFSR_66 ( );
FILL FILL_49_DFFSR_66 ( );
FILL FILL_50_DFFSR_66 ( );
FILL FILL_51_DFFSR_66 ( );
FILL FILL_0_INVX1_12 ( );
FILL FILL_1_INVX1_12 ( );
FILL FILL_2_INVX1_12 ( );
FILL FILL_3_INVX1_12 ( );
FILL FILL_0_DFFSR_90 ( );
FILL FILL_1_DFFSR_90 ( );
FILL FILL_2_DFFSR_90 ( );
FILL FILL_3_DFFSR_90 ( );
FILL FILL_4_DFFSR_90 ( );
FILL FILL_5_DFFSR_90 ( );
FILL FILL_6_DFFSR_90 ( );
FILL FILL_7_DFFSR_90 ( );
FILL FILL_8_DFFSR_90 ( );
FILL FILL_9_DFFSR_90 ( );
FILL FILL_10_DFFSR_90 ( );
FILL FILL_11_DFFSR_90 ( );
FILL FILL_12_DFFSR_90 ( );
FILL FILL_13_DFFSR_90 ( );
FILL FILL_14_DFFSR_90 ( );
FILL FILL_15_DFFSR_90 ( );
FILL FILL_16_DFFSR_90 ( );
FILL FILL_17_DFFSR_90 ( );
FILL FILL_18_DFFSR_90 ( );
FILL FILL_19_DFFSR_90 ( );
FILL FILL_20_DFFSR_90 ( );
FILL FILL_21_DFFSR_90 ( );
FILL FILL_22_DFFSR_90 ( );
FILL FILL_23_DFFSR_90 ( );
FILL FILL_24_DFFSR_90 ( );
FILL FILL_25_DFFSR_90 ( );
FILL FILL_26_DFFSR_90 ( );
FILL FILL_27_DFFSR_90 ( );
FILL FILL_28_DFFSR_90 ( );
FILL FILL_29_DFFSR_90 ( );
FILL FILL_30_DFFSR_90 ( );
FILL FILL_31_DFFSR_90 ( );
FILL FILL_32_DFFSR_90 ( );
FILL FILL_33_DFFSR_90 ( );
FILL FILL_34_DFFSR_90 ( );
FILL FILL_35_DFFSR_90 ( );
FILL FILL_36_DFFSR_90 ( );
FILL FILL_37_DFFSR_90 ( );
FILL FILL_38_DFFSR_90 ( );
FILL FILL_39_DFFSR_90 ( );
FILL FILL_40_DFFSR_90 ( );
FILL FILL_41_DFFSR_90 ( );
FILL FILL_42_DFFSR_90 ( );
FILL FILL_43_DFFSR_90 ( );
FILL FILL_44_DFFSR_90 ( );
FILL FILL_45_DFFSR_90 ( );
FILL FILL_46_DFFSR_90 ( );
FILL FILL_47_DFFSR_90 ( );
FILL FILL_48_DFFSR_90 ( );
FILL FILL_49_DFFSR_90 ( );
FILL FILL_50_DFFSR_90 ( );
FILL FILL_0_BUFX2_41 ( );
FILL FILL_1_BUFX2_41 ( );
FILL FILL_2_BUFX2_41 ( );
FILL FILL_3_BUFX2_41 ( );
FILL FILL_4_BUFX2_41 ( );
FILL FILL_5_BUFX2_41 ( );
FILL FILL_6_BUFX2_41 ( );
FILL FILL_0_DFFSR_29 ( );
FILL FILL_1_DFFSR_29 ( );
FILL FILL_2_DFFSR_29 ( );
FILL FILL_3_DFFSR_29 ( );
FILL FILL_4_DFFSR_29 ( );
FILL FILL_5_DFFSR_29 ( );
FILL FILL_6_DFFSR_29 ( );
FILL FILL_7_DFFSR_29 ( );
FILL FILL_8_DFFSR_29 ( );
FILL FILL_9_DFFSR_29 ( );
FILL FILL_10_DFFSR_29 ( );
FILL FILL_11_DFFSR_29 ( );
FILL FILL_12_DFFSR_29 ( );
FILL FILL_13_DFFSR_29 ( );
FILL FILL_14_DFFSR_29 ( );
FILL FILL_15_DFFSR_29 ( );
FILL FILL_16_DFFSR_29 ( );
FILL FILL_17_DFFSR_29 ( );
FILL FILL_18_DFFSR_29 ( );
FILL FILL_19_DFFSR_29 ( );
FILL FILL_20_DFFSR_29 ( );
FILL FILL_21_DFFSR_29 ( );
FILL FILL_22_DFFSR_29 ( );
FILL FILL_23_DFFSR_29 ( );
FILL FILL_24_DFFSR_29 ( );
FILL FILL_25_DFFSR_29 ( );
FILL FILL_26_DFFSR_29 ( );
FILL FILL_27_DFFSR_29 ( );
FILL FILL_28_DFFSR_29 ( );
FILL FILL_29_DFFSR_29 ( );
FILL FILL_30_DFFSR_29 ( );
FILL FILL_31_DFFSR_29 ( );
FILL FILL_32_DFFSR_29 ( );
FILL FILL_33_DFFSR_29 ( );
FILL FILL_34_DFFSR_29 ( );
FILL FILL_35_DFFSR_29 ( );
FILL FILL_36_DFFSR_29 ( );
FILL FILL_37_DFFSR_29 ( );
FILL FILL_38_DFFSR_29 ( );
FILL FILL_39_DFFSR_29 ( );
FILL FILL_40_DFFSR_29 ( );
FILL FILL_41_DFFSR_29 ( );
FILL FILL_42_DFFSR_29 ( );
FILL FILL_43_DFFSR_29 ( );
FILL FILL_44_DFFSR_29 ( );
FILL FILL_45_DFFSR_29 ( );
FILL FILL_46_DFFSR_29 ( );
FILL FILL_47_DFFSR_29 ( );
FILL FILL_48_DFFSR_29 ( );
FILL FILL_49_DFFSR_29 ( );
FILL FILL_50_DFFSR_29 ( );
FILL FILL_0_CLKBUF1_30 ( );
FILL FILL_1_CLKBUF1_30 ( );
FILL FILL_2_CLKBUF1_30 ( );
FILL FILL_3_CLKBUF1_30 ( );
FILL FILL_4_CLKBUF1_30 ( );
FILL FILL_5_CLKBUF1_30 ( );
FILL FILL_6_CLKBUF1_30 ( );
FILL FILL_7_CLKBUF1_30 ( );
FILL FILL_8_CLKBUF1_30 ( );
FILL FILL_9_CLKBUF1_30 ( );
FILL FILL_10_CLKBUF1_30 ( );
FILL FILL_11_CLKBUF1_30 ( );
FILL FILL_12_CLKBUF1_30 ( );
FILL FILL_13_CLKBUF1_30 ( );
FILL FILL_14_CLKBUF1_30 ( );
FILL FILL_15_CLKBUF1_30 ( );
FILL FILL_16_CLKBUF1_30 ( );
FILL FILL_17_CLKBUF1_30 ( );
FILL FILL_18_CLKBUF1_30 ( );
FILL FILL_19_CLKBUF1_30 ( );
FILL FILL_20_CLKBUF1_30 ( );
FILL FILL_0_DFFSR_133 ( );
FILL FILL_1_DFFSR_133 ( );
FILL FILL_2_DFFSR_133 ( );
FILL FILL_3_DFFSR_133 ( );
FILL FILL_4_DFFSR_133 ( );
FILL FILL_5_DFFSR_133 ( );
FILL FILL_6_DFFSR_133 ( );
FILL FILL_7_DFFSR_133 ( );
FILL FILL_8_DFFSR_133 ( );
FILL FILL_9_DFFSR_133 ( );
FILL FILL_10_DFFSR_133 ( );
FILL FILL_11_DFFSR_133 ( );
FILL FILL_12_DFFSR_133 ( );
FILL FILL_13_DFFSR_133 ( );
FILL FILL_14_DFFSR_133 ( );
FILL FILL_15_DFFSR_133 ( );
FILL FILL_16_DFFSR_133 ( );
FILL FILL_17_DFFSR_133 ( );
FILL FILL_18_DFFSR_133 ( );
FILL FILL_19_DFFSR_133 ( );
FILL FILL_20_DFFSR_133 ( );
FILL FILL_21_DFFSR_133 ( );
FILL FILL_22_DFFSR_133 ( );
FILL FILL_23_DFFSR_133 ( );
FILL FILL_24_DFFSR_133 ( );
FILL FILL_25_DFFSR_133 ( );
FILL FILL_26_DFFSR_133 ( );
FILL FILL_27_DFFSR_133 ( );
FILL FILL_28_DFFSR_133 ( );
FILL FILL_29_DFFSR_133 ( );
FILL FILL_30_DFFSR_133 ( );
FILL FILL_31_DFFSR_133 ( );
FILL FILL_32_DFFSR_133 ( );
FILL FILL_33_DFFSR_133 ( );
FILL FILL_34_DFFSR_133 ( );
FILL FILL_35_DFFSR_133 ( );
FILL FILL_36_DFFSR_133 ( );
FILL FILL_37_DFFSR_133 ( );
FILL FILL_38_DFFSR_133 ( );
FILL FILL_39_DFFSR_133 ( );
FILL FILL_40_DFFSR_133 ( );
FILL FILL_41_DFFSR_133 ( );
FILL FILL_42_DFFSR_133 ( );
FILL FILL_43_DFFSR_133 ( );
FILL FILL_44_DFFSR_133 ( );
FILL FILL_45_DFFSR_133 ( );
FILL FILL_46_DFFSR_133 ( );
FILL FILL_47_DFFSR_133 ( );
FILL FILL_48_DFFSR_133 ( );
FILL FILL_49_DFFSR_133 ( );
FILL FILL_50_DFFSR_133 ( );
FILL FILL_0_AOI22X1_16 ( );
FILL FILL_1_AOI22X1_16 ( );
FILL FILL_2_AOI22X1_16 ( );
FILL FILL_3_AOI22X1_16 ( );
FILL FILL_4_AOI22X1_16 ( );
FILL FILL_5_AOI22X1_16 ( );
FILL FILL_6_AOI22X1_16 ( );
FILL FILL_7_AOI22X1_16 ( );
FILL FILL_8_AOI22X1_16 ( );
FILL FILL_9_AOI22X1_16 ( );
FILL FILL_10_AOI22X1_16 ( );
FILL FILL_0_OAI22X1_39 ( );
FILL FILL_1_OAI22X1_39 ( );
FILL FILL_2_OAI22X1_39 ( );
FILL FILL_3_OAI22X1_39 ( );
FILL FILL_4_OAI22X1_39 ( );
FILL FILL_5_OAI22X1_39 ( );
FILL FILL_6_OAI22X1_39 ( );
FILL FILL_7_OAI22X1_39 ( );
FILL FILL_8_OAI22X1_39 ( );
FILL FILL_9_OAI22X1_39 ( );
FILL FILL_10_OAI22X1_39 ( );
FILL FILL_0_INVX1_109 ( );
FILL FILL_1_INVX1_109 ( );
FILL FILL_2_INVX1_109 ( );
FILL FILL_3_INVX1_109 ( );
FILL FILL_4_INVX1_109 ( );
FILL FILL_0_BUFX2_70 ( );
FILL FILL_1_BUFX2_70 ( );
FILL FILL_2_BUFX2_70 ( );
FILL FILL_3_BUFX2_70 ( );
FILL FILL_4_BUFX2_70 ( );
FILL FILL_5_BUFX2_70 ( );
FILL FILL_6_BUFX2_70 ( );
FILL FILL_0_INVX1_108 ( );
FILL FILL_1_INVX1_108 ( );
FILL FILL_2_INVX1_108 ( );
FILL FILL_3_INVX1_108 ( );
FILL FILL_0_DFFSR_258 ( );
FILL FILL_1_DFFSR_258 ( );
FILL FILL_2_DFFSR_258 ( );
FILL FILL_3_DFFSR_258 ( );
FILL FILL_4_DFFSR_258 ( );
FILL FILL_5_DFFSR_258 ( );
FILL FILL_6_DFFSR_258 ( );
FILL FILL_7_DFFSR_258 ( );
FILL FILL_8_DFFSR_258 ( );
FILL FILL_9_DFFSR_258 ( );
FILL FILL_10_DFFSR_258 ( );
FILL FILL_11_DFFSR_258 ( );
FILL FILL_12_DFFSR_258 ( );
FILL FILL_13_DFFSR_258 ( );
FILL FILL_14_DFFSR_258 ( );
FILL FILL_15_DFFSR_258 ( );
FILL FILL_16_DFFSR_258 ( );
FILL FILL_17_DFFSR_258 ( );
FILL FILL_18_DFFSR_258 ( );
FILL FILL_19_DFFSR_258 ( );
FILL FILL_20_DFFSR_258 ( );
FILL FILL_21_DFFSR_258 ( );
FILL FILL_22_DFFSR_258 ( );
FILL FILL_23_DFFSR_258 ( );
FILL FILL_24_DFFSR_258 ( );
FILL FILL_25_DFFSR_258 ( );
FILL FILL_26_DFFSR_258 ( );
FILL FILL_27_DFFSR_258 ( );
FILL FILL_28_DFFSR_258 ( );
FILL FILL_29_DFFSR_258 ( );
FILL FILL_30_DFFSR_258 ( );
FILL FILL_31_DFFSR_258 ( );
FILL FILL_32_DFFSR_258 ( );
FILL FILL_33_DFFSR_258 ( );
FILL FILL_34_DFFSR_258 ( );
FILL FILL_35_DFFSR_258 ( );
FILL FILL_36_DFFSR_258 ( );
FILL FILL_37_DFFSR_258 ( );
FILL FILL_38_DFFSR_258 ( );
FILL FILL_39_DFFSR_258 ( );
FILL FILL_40_DFFSR_258 ( );
FILL FILL_41_DFFSR_258 ( );
FILL FILL_42_DFFSR_258 ( );
FILL FILL_43_DFFSR_258 ( );
FILL FILL_44_DFFSR_258 ( );
FILL FILL_45_DFFSR_258 ( );
FILL FILL_46_DFFSR_258 ( );
FILL FILL_47_DFFSR_258 ( );
FILL FILL_48_DFFSR_258 ( );
FILL FILL_49_DFFSR_258 ( );
FILL FILL_50_DFFSR_258 ( );
FILL FILL_51_DFFSR_258 ( );
FILL FILL_0_INVX1_184 ( );
FILL FILL_1_INVX1_184 ( );
FILL FILL_2_INVX1_184 ( );
FILL FILL_3_INVX1_184 ( );
FILL FILL_4_INVX1_184 ( );
FILL FILL_0_OAI21X1_88 ( );
FILL FILL_1_OAI21X1_88 ( );
FILL FILL_2_OAI21X1_88 ( );
FILL FILL_3_OAI21X1_88 ( );
FILL FILL_4_OAI21X1_88 ( );
FILL FILL_5_OAI21X1_88 ( );
FILL FILL_6_OAI21X1_88 ( );
FILL FILL_7_OAI21X1_88 ( );
FILL FILL_8_OAI21X1_88 ( );
FILL FILL_0_NAND2X1_119 ( );
FILL FILL_1_NAND2X1_119 ( );
FILL FILL_2_NAND2X1_119 ( );
FILL FILL_3_NAND2X1_119 ( );
FILL FILL_4_NAND2X1_119 ( );
FILL FILL_5_NAND2X1_119 ( );
FILL FILL_6_NAND2X1_119 ( );
FILL FILL_0_DFFSR_20 ( );
FILL FILL_1_DFFSR_20 ( );
FILL FILL_2_DFFSR_20 ( );
FILL FILL_3_DFFSR_20 ( );
FILL FILL_4_DFFSR_20 ( );
FILL FILL_5_DFFSR_20 ( );
FILL FILL_6_DFFSR_20 ( );
FILL FILL_7_DFFSR_20 ( );
FILL FILL_8_DFFSR_20 ( );
FILL FILL_9_DFFSR_20 ( );
FILL FILL_10_DFFSR_20 ( );
FILL FILL_11_DFFSR_20 ( );
FILL FILL_12_DFFSR_20 ( );
FILL FILL_13_DFFSR_20 ( );
FILL FILL_14_DFFSR_20 ( );
FILL FILL_15_DFFSR_20 ( );
FILL FILL_16_DFFSR_20 ( );
FILL FILL_17_DFFSR_20 ( );
FILL FILL_18_DFFSR_20 ( );
FILL FILL_19_DFFSR_20 ( );
FILL FILL_20_DFFSR_20 ( );
FILL FILL_21_DFFSR_20 ( );
FILL FILL_22_DFFSR_20 ( );
FILL FILL_23_DFFSR_20 ( );
FILL FILL_24_DFFSR_20 ( );
FILL FILL_25_DFFSR_20 ( );
FILL FILL_26_DFFSR_20 ( );
FILL FILL_27_DFFSR_20 ( );
FILL FILL_28_DFFSR_20 ( );
FILL FILL_29_DFFSR_20 ( );
FILL FILL_30_DFFSR_20 ( );
FILL FILL_31_DFFSR_20 ( );
FILL FILL_32_DFFSR_20 ( );
FILL FILL_33_DFFSR_20 ( );
FILL FILL_34_DFFSR_20 ( );
FILL FILL_35_DFFSR_20 ( );
FILL FILL_36_DFFSR_20 ( );
FILL FILL_37_DFFSR_20 ( );
FILL FILL_38_DFFSR_20 ( );
FILL FILL_39_DFFSR_20 ( );
FILL FILL_40_DFFSR_20 ( );
FILL FILL_41_DFFSR_20 ( );
FILL FILL_42_DFFSR_20 ( );
FILL FILL_43_DFFSR_20 ( );
FILL FILL_44_DFFSR_20 ( );
FILL FILL_45_DFFSR_20 ( );
FILL FILL_46_DFFSR_20 ( );
FILL FILL_47_DFFSR_20 ( );
FILL FILL_48_DFFSR_20 ( );
FILL FILL_49_DFFSR_20 ( );
FILL FILL_50_DFFSR_20 ( );
FILL FILL_0_DFFSR_10 ( );
FILL FILL_1_DFFSR_10 ( );
FILL FILL_2_DFFSR_10 ( );
FILL FILL_3_DFFSR_10 ( );
FILL FILL_4_DFFSR_10 ( );
FILL FILL_5_DFFSR_10 ( );
FILL FILL_6_DFFSR_10 ( );
FILL FILL_7_DFFSR_10 ( );
FILL FILL_8_DFFSR_10 ( );
FILL FILL_9_DFFSR_10 ( );
FILL FILL_10_DFFSR_10 ( );
FILL FILL_11_DFFSR_10 ( );
FILL FILL_12_DFFSR_10 ( );
FILL FILL_13_DFFSR_10 ( );
FILL FILL_14_DFFSR_10 ( );
FILL FILL_15_DFFSR_10 ( );
FILL FILL_16_DFFSR_10 ( );
FILL FILL_17_DFFSR_10 ( );
FILL FILL_18_DFFSR_10 ( );
FILL FILL_19_DFFSR_10 ( );
FILL FILL_20_DFFSR_10 ( );
FILL FILL_21_DFFSR_10 ( );
FILL FILL_22_DFFSR_10 ( );
FILL FILL_23_DFFSR_10 ( );
FILL FILL_24_DFFSR_10 ( );
FILL FILL_25_DFFSR_10 ( );
FILL FILL_26_DFFSR_10 ( );
FILL FILL_27_DFFSR_10 ( );
FILL FILL_28_DFFSR_10 ( );
FILL FILL_29_DFFSR_10 ( );
FILL FILL_30_DFFSR_10 ( );
FILL FILL_31_DFFSR_10 ( );
FILL FILL_32_DFFSR_10 ( );
FILL FILL_33_DFFSR_10 ( );
FILL FILL_34_DFFSR_10 ( );
FILL FILL_35_DFFSR_10 ( );
FILL FILL_36_DFFSR_10 ( );
FILL FILL_37_DFFSR_10 ( );
FILL FILL_38_DFFSR_10 ( );
FILL FILL_39_DFFSR_10 ( );
FILL FILL_40_DFFSR_10 ( );
FILL FILL_41_DFFSR_10 ( );
FILL FILL_42_DFFSR_10 ( );
FILL FILL_43_DFFSR_10 ( );
FILL FILL_44_DFFSR_10 ( );
FILL FILL_45_DFFSR_10 ( );
FILL FILL_46_DFFSR_10 ( );
FILL FILL_47_DFFSR_10 ( );
FILL FILL_48_DFFSR_10 ( );
FILL FILL_49_DFFSR_10 ( );
FILL FILL_50_DFFSR_10 ( );
FILL FILL_0_BUFX2_71 ( );
FILL FILL_1_BUFX2_71 ( );
FILL FILL_2_BUFX2_71 ( );
FILL FILL_3_BUFX2_71 ( );
FILL FILL_4_BUFX2_71 ( );
FILL FILL_5_BUFX2_71 ( );
FILL FILL_6_BUFX2_71 ( );
FILL FILL_0_DFFSR_95 ( );
FILL FILL_1_DFFSR_95 ( );
FILL FILL_2_DFFSR_95 ( );
FILL FILL_3_DFFSR_95 ( );
FILL FILL_4_DFFSR_95 ( );
FILL FILL_5_DFFSR_95 ( );
FILL FILL_6_DFFSR_95 ( );
FILL FILL_7_DFFSR_95 ( );
FILL FILL_8_DFFSR_95 ( );
FILL FILL_9_DFFSR_95 ( );
FILL FILL_10_DFFSR_95 ( );
FILL FILL_11_DFFSR_95 ( );
FILL FILL_12_DFFSR_95 ( );
FILL FILL_13_DFFSR_95 ( );
FILL FILL_14_DFFSR_95 ( );
FILL FILL_15_DFFSR_95 ( );
FILL FILL_16_DFFSR_95 ( );
FILL FILL_17_DFFSR_95 ( );
FILL FILL_18_DFFSR_95 ( );
FILL FILL_19_DFFSR_95 ( );
FILL FILL_20_DFFSR_95 ( );
FILL FILL_21_DFFSR_95 ( );
FILL FILL_22_DFFSR_95 ( );
FILL FILL_23_DFFSR_95 ( );
FILL FILL_24_DFFSR_95 ( );
FILL FILL_25_DFFSR_95 ( );
FILL FILL_26_DFFSR_95 ( );
FILL FILL_27_DFFSR_95 ( );
FILL FILL_28_DFFSR_95 ( );
FILL FILL_29_DFFSR_95 ( );
FILL FILL_30_DFFSR_95 ( );
FILL FILL_31_DFFSR_95 ( );
FILL FILL_32_DFFSR_95 ( );
FILL FILL_33_DFFSR_95 ( );
FILL FILL_34_DFFSR_95 ( );
FILL FILL_35_DFFSR_95 ( );
FILL FILL_36_DFFSR_95 ( );
FILL FILL_37_DFFSR_95 ( );
FILL FILL_38_DFFSR_95 ( );
FILL FILL_39_DFFSR_95 ( );
FILL FILL_40_DFFSR_95 ( );
FILL FILL_41_DFFSR_95 ( );
FILL FILL_42_DFFSR_95 ( );
FILL FILL_43_DFFSR_95 ( );
FILL FILL_44_DFFSR_95 ( );
FILL FILL_45_DFFSR_95 ( );
FILL FILL_46_DFFSR_95 ( );
FILL FILL_47_DFFSR_95 ( );
FILL FILL_48_DFFSR_95 ( );
FILL FILL_49_DFFSR_95 ( );
FILL FILL_50_DFFSR_95 ( );
FILL FILL_51_DFFSR_95 ( );
FILL FILL_0_DFFSR_74 ( );
FILL FILL_1_DFFSR_74 ( );
FILL FILL_2_DFFSR_74 ( );
FILL FILL_3_DFFSR_74 ( );
FILL FILL_4_DFFSR_74 ( );
FILL FILL_5_DFFSR_74 ( );
FILL FILL_6_DFFSR_74 ( );
FILL FILL_7_DFFSR_74 ( );
FILL FILL_8_DFFSR_74 ( );
FILL FILL_9_DFFSR_74 ( );
FILL FILL_10_DFFSR_74 ( );
FILL FILL_11_DFFSR_74 ( );
FILL FILL_12_DFFSR_74 ( );
FILL FILL_13_DFFSR_74 ( );
FILL FILL_14_DFFSR_74 ( );
FILL FILL_15_DFFSR_74 ( );
FILL FILL_16_DFFSR_74 ( );
FILL FILL_17_DFFSR_74 ( );
FILL FILL_18_DFFSR_74 ( );
FILL FILL_19_DFFSR_74 ( );
FILL FILL_20_DFFSR_74 ( );
FILL FILL_21_DFFSR_74 ( );
FILL FILL_22_DFFSR_74 ( );
FILL FILL_23_DFFSR_74 ( );
FILL FILL_24_DFFSR_74 ( );
FILL FILL_25_DFFSR_74 ( );
FILL FILL_26_DFFSR_74 ( );
FILL FILL_27_DFFSR_74 ( );
FILL FILL_28_DFFSR_74 ( );
FILL FILL_29_DFFSR_74 ( );
FILL FILL_30_DFFSR_74 ( );
FILL FILL_31_DFFSR_74 ( );
FILL FILL_32_DFFSR_74 ( );
FILL FILL_33_DFFSR_74 ( );
FILL FILL_34_DFFSR_74 ( );
FILL FILL_35_DFFSR_74 ( );
FILL FILL_36_DFFSR_74 ( );
FILL FILL_37_DFFSR_74 ( );
FILL FILL_38_DFFSR_74 ( );
FILL FILL_39_DFFSR_74 ( );
FILL FILL_40_DFFSR_74 ( );
FILL FILL_41_DFFSR_74 ( );
FILL FILL_42_DFFSR_74 ( );
FILL FILL_43_DFFSR_74 ( );
FILL FILL_44_DFFSR_74 ( );
FILL FILL_45_DFFSR_74 ( );
FILL FILL_46_DFFSR_74 ( );
FILL FILL_47_DFFSR_74 ( );
FILL FILL_48_DFFSR_74 ( );
FILL FILL_49_DFFSR_74 ( );
FILL FILL_50_DFFSR_74 ( );
FILL FILL_0_CLKBUF1_35 ( );
FILL FILL_1_CLKBUF1_35 ( );
FILL FILL_2_CLKBUF1_35 ( );
FILL FILL_3_CLKBUF1_35 ( );
FILL FILL_4_CLKBUF1_35 ( );
FILL FILL_5_CLKBUF1_35 ( );
FILL FILL_6_CLKBUF1_35 ( );
FILL FILL_7_CLKBUF1_35 ( );
FILL FILL_8_CLKBUF1_35 ( );
FILL FILL_9_CLKBUF1_35 ( );
FILL FILL_10_CLKBUF1_35 ( );
FILL FILL_11_CLKBUF1_35 ( );
FILL FILL_12_CLKBUF1_35 ( );
FILL FILL_13_CLKBUF1_35 ( );
FILL FILL_14_CLKBUF1_35 ( );
FILL FILL_15_CLKBUF1_35 ( );
FILL FILL_16_CLKBUF1_35 ( );
FILL FILL_17_CLKBUF1_35 ( );
FILL FILL_18_CLKBUF1_35 ( );
FILL FILL_19_CLKBUF1_35 ( );
FILL FILL_20_CLKBUF1_35 ( );
FILL FILL_0_DFFSR_21 ( );
FILL FILL_1_DFFSR_21 ( );
FILL FILL_2_DFFSR_21 ( );
FILL FILL_3_DFFSR_21 ( );
FILL FILL_4_DFFSR_21 ( );
FILL FILL_5_DFFSR_21 ( );
FILL FILL_6_DFFSR_21 ( );
FILL FILL_7_DFFSR_21 ( );
FILL FILL_8_DFFSR_21 ( );
FILL FILL_9_DFFSR_21 ( );
FILL FILL_10_DFFSR_21 ( );
FILL FILL_11_DFFSR_21 ( );
FILL FILL_12_DFFSR_21 ( );
FILL FILL_13_DFFSR_21 ( );
FILL FILL_14_DFFSR_21 ( );
FILL FILL_15_DFFSR_21 ( );
FILL FILL_16_DFFSR_21 ( );
FILL FILL_17_DFFSR_21 ( );
FILL FILL_18_DFFSR_21 ( );
FILL FILL_19_DFFSR_21 ( );
FILL FILL_20_DFFSR_21 ( );
FILL FILL_21_DFFSR_21 ( );
FILL FILL_22_DFFSR_21 ( );
FILL FILL_23_DFFSR_21 ( );
FILL FILL_24_DFFSR_21 ( );
FILL FILL_25_DFFSR_21 ( );
FILL FILL_26_DFFSR_21 ( );
FILL FILL_27_DFFSR_21 ( );
FILL FILL_28_DFFSR_21 ( );
FILL FILL_29_DFFSR_21 ( );
FILL FILL_30_DFFSR_21 ( );
FILL FILL_31_DFFSR_21 ( );
FILL FILL_32_DFFSR_21 ( );
FILL FILL_33_DFFSR_21 ( );
FILL FILL_34_DFFSR_21 ( );
FILL FILL_35_DFFSR_21 ( );
FILL FILL_36_DFFSR_21 ( );
FILL FILL_37_DFFSR_21 ( );
FILL FILL_38_DFFSR_21 ( );
FILL FILL_39_DFFSR_21 ( );
FILL FILL_40_DFFSR_21 ( );
FILL FILL_41_DFFSR_21 ( );
FILL FILL_42_DFFSR_21 ( );
FILL FILL_43_DFFSR_21 ( );
FILL FILL_44_DFFSR_21 ( );
FILL FILL_45_DFFSR_21 ( );
FILL FILL_46_DFFSR_21 ( );
FILL FILL_47_DFFSR_21 ( );
FILL FILL_48_DFFSR_21 ( );
FILL FILL_49_DFFSR_21 ( );
FILL FILL_50_DFFSR_21 ( );
FILL FILL_51_DFFSR_21 ( );
FILL FILL_0_DFFSR_125 ( );
FILL FILL_1_DFFSR_125 ( );
FILL FILL_2_DFFSR_125 ( );
FILL FILL_3_DFFSR_125 ( );
FILL FILL_4_DFFSR_125 ( );
FILL FILL_5_DFFSR_125 ( );
FILL FILL_6_DFFSR_125 ( );
FILL FILL_7_DFFSR_125 ( );
FILL FILL_8_DFFSR_125 ( );
FILL FILL_9_DFFSR_125 ( );
FILL FILL_10_DFFSR_125 ( );
FILL FILL_11_DFFSR_125 ( );
FILL FILL_12_DFFSR_125 ( );
FILL FILL_13_DFFSR_125 ( );
FILL FILL_14_DFFSR_125 ( );
FILL FILL_15_DFFSR_125 ( );
FILL FILL_16_DFFSR_125 ( );
FILL FILL_17_DFFSR_125 ( );
FILL FILL_18_DFFSR_125 ( );
FILL FILL_19_DFFSR_125 ( );
FILL FILL_20_DFFSR_125 ( );
FILL FILL_21_DFFSR_125 ( );
FILL FILL_22_DFFSR_125 ( );
FILL FILL_23_DFFSR_125 ( );
FILL FILL_24_DFFSR_125 ( );
FILL FILL_25_DFFSR_125 ( );
FILL FILL_26_DFFSR_125 ( );
FILL FILL_27_DFFSR_125 ( );
FILL FILL_28_DFFSR_125 ( );
FILL FILL_29_DFFSR_125 ( );
FILL FILL_30_DFFSR_125 ( );
FILL FILL_31_DFFSR_125 ( );
FILL FILL_32_DFFSR_125 ( );
FILL FILL_33_DFFSR_125 ( );
FILL FILL_34_DFFSR_125 ( );
FILL FILL_35_DFFSR_125 ( );
FILL FILL_36_DFFSR_125 ( );
FILL FILL_37_DFFSR_125 ( );
FILL FILL_38_DFFSR_125 ( );
FILL FILL_39_DFFSR_125 ( );
FILL FILL_40_DFFSR_125 ( );
FILL FILL_41_DFFSR_125 ( );
FILL FILL_42_DFFSR_125 ( );
FILL FILL_43_DFFSR_125 ( );
FILL FILL_44_DFFSR_125 ( );
FILL FILL_45_DFFSR_125 ( );
FILL FILL_46_DFFSR_125 ( );
FILL FILL_47_DFFSR_125 ( );
FILL FILL_48_DFFSR_125 ( );
FILL FILL_49_DFFSR_125 ( );
FILL FILL_50_DFFSR_125 ( );
FILL FILL_0_NAND3X1_77 ( );
FILL FILL_1_NAND3X1_77 ( );
FILL FILL_2_NAND3X1_77 ( );
FILL FILL_3_NAND3X1_77 ( );
FILL FILL_4_NAND3X1_77 ( );
FILL FILL_5_NAND3X1_77 ( );
FILL FILL_6_NAND3X1_77 ( );
FILL FILL_7_NAND3X1_77 ( );
FILL FILL_8_NAND3X1_77 ( );
FILL FILL_0_INVX1_116 ( );
FILL FILL_1_INVX1_116 ( );
FILL FILL_2_INVX1_116 ( );
FILL FILL_3_INVX1_116 ( );
FILL FILL_4_INVX1_116 ( );
FILL FILL_0_DFFSR_5 ( );
FILL FILL_1_DFFSR_5 ( );
FILL FILL_2_DFFSR_5 ( );
FILL FILL_3_DFFSR_5 ( );
FILL FILL_4_DFFSR_5 ( );
FILL FILL_5_DFFSR_5 ( );
FILL FILL_6_DFFSR_5 ( );
FILL FILL_7_DFFSR_5 ( );
FILL FILL_8_DFFSR_5 ( );
FILL FILL_9_DFFSR_5 ( );
FILL FILL_10_DFFSR_5 ( );
FILL FILL_11_DFFSR_5 ( );
FILL FILL_12_DFFSR_5 ( );
FILL FILL_13_DFFSR_5 ( );
FILL FILL_14_DFFSR_5 ( );
FILL FILL_15_DFFSR_5 ( );
FILL FILL_16_DFFSR_5 ( );
FILL FILL_17_DFFSR_5 ( );
FILL FILL_18_DFFSR_5 ( );
FILL FILL_19_DFFSR_5 ( );
FILL FILL_20_DFFSR_5 ( );
FILL FILL_21_DFFSR_5 ( );
FILL FILL_22_DFFSR_5 ( );
FILL FILL_23_DFFSR_5 ( );
FILL FILL_24_DFFSR_5 ( );
FILL FILL_25_DFFSR_5 ( );
FILL FILL_26_DFFSR_5 ( );
FILL FILL_27_DFFSR_5 ( );
FILL FILL_28_DFFSR_5 ( );
FILL FILL_29_DFFSR_5 ( );
FILL FILL_30_DFFSR_5 ( );
FILL FILL_31_DFFSR_5 ( );
FILL FILL_32_DFFSR_5 ( );
FILL FILL_33_DFFSR_5 ( );
FILL FILL_34_DFFSR_5 ( );
FILL FILL_35_DFFSR_5 ( );
FILL FILL_36_DFFSR_5 ( );
FILL FILL_37_DFFSR_5 ( );
FILL FILL_38_DFFSR_5 ( );
FILL FILL_39_DFFSR_5 ( );
FILL FILL_40_DFFSR_5 ( );
FILL FILL_41_DFFSR_5 ( );
FILL FILL_42_DFFSR_5 ( );
FILL FILL_43_DFFSR_5 ( );
FILL FILL_44_DFFSR_5 ( );
FILL FILL_45_DFFSR_5 ( );
FILL FILL_46_DFFSR_5 ( );
FILL FILL_47_DFFSR_5 ( );
FILL FILL_48_DFFSR_5 ( );
FILL FILL_49_DFFSR_5 ( );
FILL FILL_50_DFFSR_5 ( );
FILL FILL_0_0_0 ( );
FILL FILL_0_0_1 ( );
FILL FILL_0_0_2 ( );
FILL FILL_0_1_0 ( );
FILL FILL_0_1_1 ( );
FILL FILL_0_1_2 ( );
FILL FILL_0_2_0 ( );
FILL FILL_0_2_1 ( );
FILL FILL_0_2_2 ( );
FILL FILL_0_3_0 ( );
FILL FILL_0_3_1 ( );
FILL FILL_0_3_2 ( );
FILL FILL_0_4_0 ( );
FILL FILL_0_4_1 ( );
FILL FILL_0_4_2 ( );
FILL FILL_0_5_0 ( );
FILL FILL_0_5_1 ( );
FILL FILL_0_5_2 ( );
FILL FILL_0_6_0 ( );
FILL FILL_0_6_1 ( );
FILL FILL_0_6_2 ( );
FILL FILL_1_1 ( );
FILL FILL_1_2 ( );
FILL FILL_1_3 ( );
FILL FILL_1_4 ( );
FILL FILL_1_5 ( );
FILL FILL_1_6 ( );
FILL FILL_1_7 ( );
FILL FILL_1_0_0 ( );
FILL FILL_1_0_1 ( );
FILL FILL_1_0_2 ( );
FILL FILL_1_1_0 ( );
FILL FILL_1_1_1 ( );
FILL FILL_1_1_2 ( );
FILL FILL_1_2_0 ( );
FILL FILL_1_2_1 ( );
FILL FILL_1_2_2 ( );
FILL FILL_1_3_0 ( );
FILL FILL_1_3_1 ( );
FILL FILL_1_3_2 ( );
FILL FILL_1_4_0 ( );
FILL FILL_1_4_1 ( );
FILL FILL_1_4_2 ( );
FILL FILL_1_5_0 ( );
FILL FILL_1_5_1 ( );
FILL FILL_1_5_2 ( );
FILL FILL_1_6_0 ( );
FILL FILL_1_6_1 ( );
FILL FILL_1_6_2 ( );
FILL FILL_2_1 ( );
FILL FILL_2_0_0 ( );
FILL FILL_2_0_1 ( );
FILL FILL_2_0_2 ( );
FILL FILL_2_1_0 ( );
FILL FILL_2_1_1 ( );
FILL FILL_2_1_2 ( );
FILL FILL_2_2_0 ( );
FILL FILL_2_2_1 ( );
FILL FILL_2_2_2 ( );
FILL FILL_2_3_0 ( );
FILL FILL_2_3_1 ( );
FILL FILL_2_3_2 ( );
FILL FILL_2_4_0 ( );
FILL FILL_2_4_1 ( );
FILL FILL_2_4_2 ( );
FILL FILL_2_5_0 ( );
FILL FILL_2_5_1 ( );
FILL FILL_2_5_2 ( );
FILL FILL_2_6_0 ( );
FILL FILL_2_6_1 ( );
FILL FILL_2_6_2 ( );
FILL FILL_3_1 ( );
FILL FILL_3_2 ( );
FILL FILL_3_3 ( );
FILL FILL_3_4 ( );
FILL FILL_3_0_0 ( );
FILL FILL_3_0_1 ( );
FILL FILL_3_0_2 ( );
FILL FILL_3_1_0 ( );
FILL FILL_3_1_1 ( );
FILL FILL_3_1_2 ( );
FILL FILL_3_2_0 ( );
FILL FILL_3_2_1 ( );
FILL FILL_3_2_2 ( );
FILL FILL_3_3_0 ( );
FILL FILL_3_3_1 ( );
FILL FILL_3_3_2 ( );
FILL FILL_3_4_0 ( );
FILL FILL_3_4_1 ( );
FILL FILL_3_4_2 ( );
FILL FILL_3_5_0 ( );
FILL FILL_3_5_1 ( );
FILL FILL_3_5_2 ( );
FILL FILL_3_6_0 ( );
FILL FILL_3_6_1 ( );
FILL FILL_3_6_2 ( );
FILL FILL_4_1 ( );
FILL FILL_4_0_0 ( );
FILL FILL_4_0_1 ( );
FILL FILL_4_0_2 ( );
FILL FILL_4_1_0 ( );
FILL FILL_4_1_1 ( );
FILL FILL_4_1_2 ( );
FILL FILL_4_2_0 ( );
FILL FILL_4_2_1 ( );
FILL FILL_4_2_2 ( );
FILL FILL_4_3_0 ( );
FILL FILL_4_3_1 ( );
FILL FILL_4_3_2 ( );
FILL FILL_4_4_0 ( );
FILL FILL_4_4_1 ( );
FILL FILL_4_4_2 ( );
FILL FILL_4_5_0 ( );
FILL FILL_4_5_1 ( );
FILL FILL_4_5_2 ( );
FILL FILL_4_6_0 ( );
FILL FILL_4_6_1 ( );
FILL FILL_4_6_2 ( );
FILL FILL_5_1 ( );
FILL FILL_5_2 ( );
FILL FILL_5_3 ( );
FILL FILL_5_4 ( );
FILL FILL_5_5 ( );
FILL FILL_5_6 ( );
FILL FILL_5_7 ( );
FILL FILL_5_8 ( );
FILL FILL_5_9 ( );
FILL FILL_5_10 ( );
FILL FILL_5_0_0 ( );
FILL FILL_5_0_1 ( );
FILL FILL_5_0_2 ( );
FILL FILL_5_1_0 ( );
FILL FILL_5_1_1 ( );
FILL FILL_5_1_2 ( );
FILL FILL_5_2_0 ( );
FILL FILL_5_2_1 ( );
FILL FILL_5_2_2 ( );
FILL FILL_5_3_0 ( );
FILL FILL_5_3_1 ( );
FILL FILL_5_3_2 ( );
FILL FILL_5_4_0 ( );
FILL FILL_5_4_1 ( );
FILL FILL_5_4_2 ( );
FILL FILL_5_5_0 ( );
FILL FILL_5_5_1 ( );
FILL FILL_5_5_2 ( );
FILL FILL_5_6_0 ( );
FILL FILL_5_6_1 ( );
FILL FILL_5_6_2 ( );
FILL FILL_6_1 ( );
FILL FILL_6_0_0 ( );
FILL FILL_6_0_1 ( );
FILL FILL_6_0_2 ( );
FILL FILL_6_1_0 ( );
FILL FILL_6_1_1 ( );
FILL FILL_6_1_2 ( );
FILL FILL_6_2_0 ( );
FILL FILL_6_2_1 ( );
FILL FILL_6_2_2 ( );
FILL FILL_6_3_0 ( );
FILL FILL_6_3_1 ( );
FILL FILL_6_3_2 ( );
FILL FILL_6_4_0 ( );
FILL FILL_6_4_1 ( );
FILL FILL_6_4_2 ( );
FILL FILL_6_5_0 ( );
FILL FILL_6_5_1 ( );
FILL FILL_6_5_2 ( );
FILL FILL_6_6_0 ( );
FILL FILL_6_6_1 ( );
FILL FILL_6_6_2 ( );
FILL FILL_7_1 ( );
FILL FILL_7_2 ( );
FILL FILL_7_3 ( );
FILL FILL_7_4 ( );
FILL FILL_7_5 ( );
FILL FILL_7_6 ( );
FILL FILL_7_7 ( );
FILL FILL_7_8 ( );
FILL FILL_7_9 ( );
FILL FILL_7_10 ( );
FILL FILL_7_0_0 ( );
FILL FILL_7_0_1 ( );
FILL FILL_7_0_2 ( );
FILL FILL_7_1_0 ( );
FILL FILL_7_1_1 ( );
FILL FILL_7_1_2 ( );
FILL FILL_7_2_0 ( );
FILL FILL_7_2_1 ( );
FILL FILL_7_2_2 ( );
FILL FILL_7_3_0 ( );
FILL FILL_7_3_1 ( );
FILL FILL_7_3_2 ( );
FILL FILL_7_4_0 ( );
FILL FILL_7_4_1 ( );
FILL FILL_7_4_2 ( );
FILL FILL_7_5_0 ( );
FILL FILL_7_5_1 ( );
FILL FILL_7_5_2 ( );
FILL FILL_7_6_0 ( );
FILL FILL_7_6_1 ( );
FILL FILL_7_6_2 ( );
FILL FILL_8_1 ( );
FILL FILL_8_2 ( );
FILL FILL_8_3 ( );
FILL FILL_8_4 ( );
FILL FILL_8_5 ( );
FILL FILL_8_6 ( );
FILL FILL_8_7 ( );
FILL FILL_8_8 ( );
FILL FILL_8_0_0 ( );
FILL FILL_8_0_1 ( );
FILL FILL_8_0_2 ( );
FILL FILL_8_1_0 ( );
FILL FILL_8_1_1 ( );
FILL FILL_8_1_2 ( );
FILL FILL_8_2_0 ( );
FILL FILL_8_2_1 ( );
FILL FILL_8_2_2 ( );
FILL FILL_8_3_0 ( );
FILL FILL_8_3_1 ( );
FILL FILL_8_3_2 ( );
FILL FILL_8_4_0 ( );
FILL FILL_8_4_1 ( );
FILL FILL_8_4_2 ( );
FILL FILL_8_5_0 ( );
FILL FILL_8_5_1 ( );
FILL FILL_8_5_2 ( );
FILL FILL_8_6_0 ( );
FILL FILL_8_6_1 ( );
FILL FILL_8_6_2 ( );
FILL FILL_9_1 ( );
FILL FILL_9_2 ( );
FILL FILL_9_3 ( );
FILL FILL_9_4 ( );
FILL FILL_9_5 ( );
FILL FILL_9_6 ( );
FILL FILL_9_0_0 ( );
FILL FILL_9_0_1 ( );
FILL FILL_9_0_2 ( );
FILL FILL_9_1_0 ( );
FILL FILL_9_1_1 ( );
FILL FILL_9_1_2 ( );
FILL FILL_9_2_0 ( );
FILL FILL_9_2_1 ( );
FILL FILL_9_2_2 ( );
FILL FILL_9_3_0 ( );
FILL FILL_9_3_1 ( );
FILL FILL_9_3_2 ( );
FILL FILL_9_4_0 ( );
FILL FILL_9_4_1 ( );
FILL FILL_9_4_2 ( );
FILL FILL_9_5_0 ( );
FILL FILL_9_5_1 ( );
FILL FILL_9_5_2 ( );
FILL FILL_9_6_0 ( );
FILL FILL_9_6_1 ( );
FILL FILL_9_6_2 ( );
FILL FILL_10_1 ( );
FILL FILL_10_2 ( );
FILL FILL_10_3 ( );
FILL FILL_10_4 ( );
FILL FILL_10_5 ( );
FILL FILL_10_6 ( );
FILL FILL_10_0_0 ( );
FILL FILL_10_0_1 ( );
FILL FILL_10_0_2 ( );
FILL FILL_10_1_0 ( );
FILL FILL_10_1_1 ( );
FILL FILL_10_1_2 ( );
FILL FILL_10_2_0 ( );
FILL FILL_10_2_1 ( );
FILL FILL_10_2_2 ( );
FILL FILL_10_3_0 ( );
FILL FILL_10_3_1 ( );
FILL FILL_10_3_2 ( );
FILL FILL_10_4_0 ( );
FILL FILL_10_4_1 ( );
FILL FILL_10_4_2 ( );
FILL FILL_10_5_0 ( );
FILL FILL_10_5_1 ( );
FILL FILL_10_5_2 ( );
FILL FILL_10_6_0 ( );
FILL FILL_10_6_1 ( );
FILL FILL_10_6_2 ( );
FILL FILL_11_1 ( );
FILL FILL_11_2 ( );
FILL FILL_11_3 ( );
FILL FILL_11_4 ( );
FILL FILL_11_5 ( );
FILL FILL_11_6 ( );
FILL FILL_11_7 ( );
FILL FILL_11_0_0 ( );
FILL FILL_11_0_1 ( );
FILL FILL_11_0_2 ( );
FILL FILL_11_1_0 ( );
FILL FILL_11_1_1 ( );
FILL FILL_11_1_2 ( );
FILL FILL_11_2_0 ( );
FILL FILL_11_2_1 ( );
FILL FILL_11_2_2 ( );
FILL FILL_11_3_0 ( );
FILL FILL_11_3_1 ( );
FILL FILL_11_3_2 ( );
FILL FILL_11_4_0 ( );
FILL FILL_11_4_1 ( );
FILL FILL_11_4_2 ( );
FILL FILL_11_5_0 ( );
FILL FILL_11_5_1 ( );
FILL FILL_11_5_2 ( );
FILL FILL_11_6_0 ( );
FILL FILL_11_6_1 ( );
FILL FILL_11_6_2 ( );
FILL FILL_12_1 ( );
FILL FILL_12_2 ( );
FILL FILL_12_3 ( );
FILL FILL_12_0_0 ( );
FILL FILL_12_0_1 ( );
FILL FILL_12_0_2 ( );
FILL FILL_12_1_0 ( );
FILL FILL_12_1_1 ( );
FILL FILL_12_1_2 ( );
FILL FILL_12_2_0 ( );
FILL FILL_12_2_1 ( );
FILL FILL_12_2_2 ( );
FILL FILL_12_3_0 ( );
FILL FILL_12_3_1 ( );
FILL FILL_12_3_2 ( );
FILL FILL_12_4_0 ( );
FILL FILL_12_4_1 ( );
FILL FILL_12_4_2 ( );
FILL FILL_12_5_0 ( );
FILL FILL_12_5_1 ( );
FILL FILL_12_5_2 ( );
FILL FILL_12_6_0 ( );
FILL FILL_12_6_1 ( );
FILL FILL_12_6_2 ( );
FILL FILL_13_1 ( );
FILL FILL_13_2 ( );
FILL FILL_13_0_0 ( );
FILL FILL_13_0_1 ( );
FILL FILL_13_0_2 ( );
FILL FILL_13_1_0 ( );
FILL FILL_13_1_1 ( );
FILL FILL_13_1_2 ( );
FILL FILL_13_2_0 ( );
FILL FILL_13_2_1 ( );
FILL FILL_13_2_2 ( );
FILL FILL_13_3_0 ( );
FILL FILL_13_3_1 ( );
FILL FILL_13_3_2 ( );
FILL FILL_13_4_0 ( );
FILL FILL_13_4_1 ( );
FILL FILL_13_4_2 ( );
FILL FILL_13_5_0 ( );
FILL FILL_13_5_1 ( );
FILL FILL_13_5_2 ( );
FILL FILL_13_6_0 ( );
FILL FILL_13_6_1 ( );
FILL FILL_13_6_2 ( );
FILL FILL_14_1 ( );
FILL FILL_14_2 ( );
FILL FILL_14_3 ( );
FILL FILL_14_4 ( );
FILL FILL_14_5 ( );
FILL FILL_14_0_0 ( );
FILL FILL_14_0_1 ( );
FILL FILL_14_0_2 ( );
FILL FILL_14_1_0 ( );
FILL FILL_14_1_1 ( );
FILL FILL_14_1_2 ( );
FILL FILL_14_2_0 ( );
FILL FILL_14_2_1 ( );
FILL FILL_14_2_2 ( );
FILL FILL_14_3_0 ( );
FILL FILL_14_3_1 ( );
FILL FILL_14_3_2 ( );
FILL FILL_14_4_0 ( );
FILL FILL_14_4_1 ( );
FILL FILL_14_4_2 ( );
FILL FILL_14_5_0 ( );
FILL FILL_14_5_1 ( );
FILL FILL_14_5_2 ( );
FILL FILL_14_6_0 ( );
FILL FILL_14_6_1 ( );
FILL FILL_14_6_2 ( );
FILL FILL_15_1 ( );
FILL FILL_15_2 ( );
FILL FILL_15_3 ( );
FILL FILL_15_4 ( );
FILL FILL_15_5 ( );
FILL FILL_15_0_0 ( );
FILL FILL_15_0_1 ( );
FILL FILL_15_0_2 ( );
FILL FILL_15_1_0 ( );
FILL FILL_15_1_1 ( );
FILL FILL_15_1_2 ( );
FILL FILL_15_2_0 ( );
FILL FILL_15_2_1 ( );
FILL FILL_15_2_2 ( );
FILL FILL_15_3_0 ( );
FILL FILL_15_3_1 ( );
FILL FILL_15_3_2 ( );
FILL FILL_15_4_0 ( );
FILL FILL_15_4_1 ( );
FILL FILL_15_4_2 ( );
FILL FILL_15_5_0 ( );
FILL FILL_15_5_1 ( );
FILL FILL_15_5_2 ( );
FILL FILL_15_6_0 ( );
FILL FILL_15_6_1 ( );
FILL FILL_15_6_2 ( );
FILL FILL_16_1 ( );
FILL FILL_16_2 ( );
FILL FILL_16_3 ( );
FILL FILL_16_4 ( );
FILL FILL_16_0_0 ( );
FILL FILL_16_0_1 ( );
FILL FILL_16_0_2 ( );
FILL FILL_16_1_0 ( );
FILL FILL_16_1_1 ( );
FILL FILL_16_1_2 ( );
FILL FILL_16_2_0 ( );
FILL FILL_16_2_1 ( );
FILL FILL_16_2_2 ( );
FILL FILL_16_3_0 ( );
FILL FILL_16_3_1 ( );
FILL FILL_16_3_2 ( );
FILL FILL_16_4_0 ( );
FILL FILL_16_4_1 ( );
FILL FILL_16_4_2 ( );
FILL FILL_16_5_0 ( );
FILL FILL_16_5_1 ( );
FILL FILL_16_5_2 ( );
FILL FILL_16_6_0 ( );
FILL FILL_16_6_1 ( );
FILL FILL_16_6_2 ( );
FILL FILL_17_1 ( );
FILL FILL_17_2 ( );
FILL FILL_17_3 ( );
FILL FILL_17_4 ( );
FILL FILL_17_5 ( );
FILL FILL_17_6 ( );
FILL FILL_17_0_0 ( );
FILL FILL_17_0_1 ( );
FILL FILL_17_0_2 ( );
FILL FILL_17_1_0 ( );
FILL FILL_17_1_1 ( );
FILL FILL_17_1_2 ( );
FILL FILL_17_2_0 ( );
FILL FILL_17_2_1 ( );
FILL FILL_17_2_2 ( );
FILL FILL_17_3_0 ( );
FILL FILL_17_3_1 ( );
FILL FILL_17_3_2 ( );
FILL FILL_17_4_0 ( );
FILL FILL_17_4_1 ( );
FILL FILL_17_4_2 ( );
FILL FILL_17_5_0 ( );
FILL FILL_17_5_1 ( );
FILL FILL_17_5_2 ( );
FILL FILL_17_6_0 ( );
FILL FILL_17_6_1 ( );
FILL FILL_17_6_2 ( );
FILL FILL_18_1 ( );
FILL FILL_18_2 ( );
FILL FILL_18_3 ( );
FILL FILL_18_4 ( );
FILL FILL_18_5 ( );
FILL FILL_18_6 ( );
FILL FILL_18_0_0 ( );
FILL FILL_18_0_1 ( );
FILL FILL_18_0_2 ( );
FILL FILL_18_1_0 ( );
FILL FILL_18_1_1 ( );
FILL FILL_18_1_2 ( );
FILL FILL_18_2_0 ( );
FILL FILL_18_2_1 ( );
FILL FILL_18_2_2 ( );
FILL FILL_18_3_0 ( );
FILL FILL_18_3_1 ( );
FILL FILL_18_3_2 ( );
FILL FILL_18_4_0 ( );
FILL FILL_18_4_1 ( );
FILL FILL_18_4_2 ( );
FILL FILL_18_5_0 ( );
FILL FILL_18_5_1 ( );
FILL FILL_18_5_2 ( );
FILL FILL_18_6_0 ( );
FILL FILL_18_6_1 ( );
FILL FILL_18_6_2 ( );
FILL FILL_19_1 ( );
FILL FILL_19_2 ( );
FILL FILL_19_3 ( );
FILL FILL_19_4 ( );
FILL FILL_19_5 ( );
FILL FILL_19_6 ( );
FILL FILL_19_7 ( );
FILL FILL_19_8 ( );
FILL FILL_19_9 ( );
FILL FILL_19_0_0 ( );
FILL FILL_19_0_1 ( );
FILL FILL_19_0_2 ( );
FILL FILL_19_1_0 ( );
FILL FILL_19_1_1 ( );
FILL FILL_19_1_2 ( );
FILL FILL_19_2_0 ( );
FILL FILL_19_2_1 ( );
FILL FILL_19_2_2 ( );
FILL FILL_19_3_0 ( );
FILL FILL_19_3_1 ( );
FILL FILL_19_3_2 ( );
FILL FILL_19_4_0 ( );
FILL FILL_19_4_1 ( );
FILL FILL_19_4_2 ( );
FILL FILL_19_5_0 ( );
FILL FILL_19_5_1 ( );
FILL FILL_19_5_2 ( );
FILL FILL_19_6_0 ( );
FILL FILL_19_6_1 ( );
FILL FILL_19_6_2 ( );
FILL FILL_20_1 ( );
FILL FILL_20_2 ( );
FILL FILL_20_3 ( );
FILL FILL_20_4 ( );
FILL FILL_20_5 ( );
FILL FILL_20_6 ( );
FILL FILL_20_0_0 ( );
FILL FILL_20_0_1 ( );
FILL FILL_20_0_2 ( );
FILL FILL_20_1_0 ( );
FILL FILL_20_1_1 ( );
FILL FILL_20_1_2 ( );
FILL FILL_20_2_0 ( );
FILL FILL_20_2_1 ( );
FILL FILL_20_2_2 ( );
FILL FILL_20_3_0 ( );
FILL FILL_20_3_1 ( );
FILL FILL_20_3_2 ( );
FILL FILL_20_4_0 ( );
FILL FILL_20_4_1 ( );
FILL FILL_20_4_2 ( );
FILL FILL_20_5_0 ( );
FILL FILL_20_5_1 ( );
FILL FILL_20_5_2 ( );
FILL FILL_20_6_0 ( );
FILL FILL_20_6_1 ( );
FILL FILL_20_6_2 ( );
FILL FILL_21_0_0 ( );
FILL FILL_21_0_1 ( );
FILL FILL_21_0_2 ( );
FILL FILL_21_1_0 ( );
FILL FILL_21_1_1 ( );
FILL FILL_21_1_2 ( );
FILL FILL_21_2_0 ( );
FILL FILL_21_2_1 ( );
FILL FILL_21_2_2 ( );
FILL FILL_21_3_0 ( );
FILL FILL_21_3_1 ( );
FILL FILL_21_3_2 ( );
FILL FILL_21_4_0 ( );
FILL FILL_21_4_1 ( );
FILL FILL_21_4_2 ( );
FILL FILL_21_5_0 ( );
FILL FILL_21_5_1 ( );
FILL FILL_21_5_2 ( );
FILL FILL_21_6_0 ( );
FILL FILL_21_6_1 ( );
FILL FILL_21_6_2 ( );
FILL FILL_22_1 ( );
FILL FILL_22_2 ( );
FILL FILL_22_3 ( );
FILL FILL_22_4 ( );
FILL FILL_22_5 ( );
FILL FILL_22_6 ( );
FILL FILL_22_0_0 ( );
FILL FILL_22_0_1 ( );
FILL FILL_22_0_2 ( );
FILL FILL_22_1_0 ( );
FILL FILL_22_1_1 ( );
FILL FILL_22_1_2 ( );
FILL FILL_22_2_0 ( );
FILL FILL_22_2_1 ( );
FILL FILL_22_2_2 ( );
FILL FILL_22_3_0 ( );
FILL FILL_22_3_1 ( );
FILL FILL_22_3_2 ( );
FILL FILL_22_4_0 ( );
FILL FILL_22_4_1 ( );
FILL FILL_22_4_2 ( );
FILL FILL_22_5_0 ( );
FILL FILL_22_5_1 ( );
FILL FILL_22_5_2 ( );
FILL FILL_22_6_0 ( );
FILL FILL_22_6_1 ( );
FILL FILL_22_6_2 ( );
FILL FILL_23_0_0 ( );
FILL FILL_23_0_1 ( );
FILL FILL_23_0_2 ( );
FILL FILL_23_1_0 ( );
FILL FILL_23_1_1 ( );
FILL FILL_23_1_2 ( );
FILL FILL_23_2_0 ( );
FILL FILL_23_2_1 ( );
FILL FILL_23_2_2 ( );
FILL FILL_23_3_0 ( );
FILL FILL_23_3_1 ( );
FILL FILL_23_3_2 ( );
FILL FILL_23_4_0 ( );
FILL FILL_23_4_1 ( );
FILL FILL_23_4_2 ( );
FILL FILL_23_5_0 ( );
FILL FILL_23_5_1 ( );
FILL FILL_23_5_2 ( );
FILL FILL_23_6_0 ( );
FILL FILL_23_6_1 ( );
FILL FILL_23_6_2 ( );
FILL FILL_24_1 ( );
FILL FILL_24_2 ( );
FILL FILL_24_3 ( );
FILL FILL_24_4 ( );
FILL FILL_24_5 ( );
FILL FILL_24_6 ( );
FILL FILL_24_7 ( );
FILL FILL_24_8 ( );
FILL FILL_24_9 ( );
FILL FILL_24_0_0 ( );
FILL FILL_24_0_1 ( );
FILL FILL_24_0_2 ( );
FILL FILL_24_1_0 ( );
FILL FILL_24_1_1 ( );
FILL FILL_24_1_2 ( );
FILL FILL_24_2_0 ( );
FILL FILL_24_2_1 ( );
FILL FILL_24_2_2 ( );
FILL FILL_24_3_0 ( );
FILL FILL_24_3_1 ( );
FILL FILL_24_3_2 ( );
FILL FILL_24_4_0 ( );
FILL FILL_24_4_1 ( );
FILL FILL_24_4_2 ( );
FILL FILL_24_5_0 ( );
FILL FILL_24_5_1 ( );
FILL FILL_24_5_2 ( );
FILL FILL_24_6_0 ( );
FILL FILL_24_6_1 ( );
FILL FILL_24_6_2 ( );
FILL FILL_25_0_0 ( );
FILL FILL_25_0_1 ( );
FILL FILL_25_0_2 ( );
FILL FILL_25_1_0 ( );
FILL FILL_25_1_1 ( );
FILL FILL_25_1_2 ( );
FILL FILL_25_2_0 ( );
FILL FILL_25_2_1 ( );
FILL FILL_25_2_2 ( );
FILL FILL_25_3_0 ( );
FILL FILL_25_3_1 ( );
FILL FILL_25_3_2 ( );
FILL FILL_25_4_0 ( );
FILL FILL_25_4_1 ( );
FILL FILL_25_4_2 ( );
FILL FILL_25_5_0 ( );
FILL FILL_25_5_1 ( );
FILL FILL_25_5_2 ( );
FILL FILL_25_6_0 ( );
FILL FILL_25_6_1 ( );
FILL FILL_25_6_2 ( );
FILL FILL_26_1 ( );
FILL FILL_26_2 ( );
FILL FILL_26_0_0 ( );
FILL FILL_26_0_1 ( );
FILL FILL_26_0_2 ( );
FILL FILL_26_1_0 ( );
FILL FILL_26_1_1 ( );
FILL FILL_26_1_2 ( );
FILL FILL_26_2_0 ( );
FILL FILL_26_2_1 ( );
FILL FILL_26_2_2 ( );
FILL FILL_26_3_0 ( );
FILL FILL_26_3_1 ( );
FILL FILL_26_3_2 ( );
FILL FILL_26_4_0 ( );
FILL FILL_26_4_1 ( );
FILL FILL_26_4_2 ( );
FILL FILL_26_5_0 ( );
FILL FILL_26_5_1 ( );
FILL FILL_26_5_2 ( );
FILL FILL_26_6_0 ( );
FILL FILL_26_6_1 ( );
FILL FILL_26_6_2 ( );
FILL FILL_27_1 ( );
FILL FILL_27_0_0 ( );
FILL FILL_27_0_1 ( );
FILL FILL_27_0_2 ( );
FILL FILL_27_1_0 ( );
FILL FILL_27_1_1 ( );
FILL FILL_27_1_2 ( );
FILL FILL_27_2_0 ( );
FILL FILL_27_2_1 ( );
FILL FILL_27_2_2 ( );
FILL FILL_27_3_0 ( );
FILL FILL_27_3_1 ( );
FILL FILL_27_3_2 ( );
FILL FILL_27_4_0 ( );
FILL FILL_27_4_1 ( );
FILL FILL_27_4_2 ( );
FILL FILL_27_5_0 ( );
FILL FILL_27_5_1 ( );
FILL FILL_27_5_2 ( );
FILL FILL_27_6_0 ( );
FILL FILL_27_6_1 ( );
FILL FILL_27_6_2 ( );
FILL FILL_28_1 ( );
FILL FILL_28_2 ( );
FILL FILL_28_0_0 ( );
FILL FILL_28_0_1 ( );
FILL FILL_28_0_2 ( );
FILL FILL_28_1_0 ( );
FILL FILL_28_1_1 ( );
FILL FILL_28_1_2 ( );
FILL FILL_28_2_0 ( );
FILL FILL_28_2_1 ( );
FILL FILL_28_2_2 ( );
FILL FILL_28_3_0 ( );
FILL FILL_28_3_1 ( );
FILL FILL_28_3_2 ( );
FILL FILL_28_4_0 ( );
FILL FILL_28_4_1 ( );
FILL FILL_28_4_2 ( );
FILL FILL_28_5_0 ( );
FILL FILL_28_5_1 ( );
FILL FILL_28_5_2 ( );
FILL FILL_28_6_0 ( );
FILL FILL_28_6_1 ( );
FILL FILL_28_6_2 ( );
FILL FILL_29_0_0 ( );
FILL FILL_29_0_1 ( );
FILL FILL_29_0_2 ( );
FILL FILL_29_1_0 ( );
FILL FILL_29_1_1 ( );
FILL FILL_29_1_2 ( );
FILL FILL_29_2_0 ( );
FILL FILL_29_2_1 ( );
FILL FILL_29_2_2 ( );
FILL FILL_29_3_0 ( );
FILL FILL_29_3_1 ( );
FILL FILL_29_3_2 ( );
FILL FILL_29_4_0 ( );
FILL FILL_29_4_1 ( );
FILL FILL_29_4_2 ( );
FILL FILL_29_5_0 ( );
FILL FILL_29_5_1 ( );
FILL FILL_29_5_2 ( );
FILL FILL_29_6_0 ( );
FILL FILL_29_6_1 ( );
FILL FILL_29_6_2 ( );
FILL FILL_30_1 ( );
FILL FILL_30_2 ( );
FILL FILL_30_3 ( );
FILL FILL_30_4 ( );
FILL FILL_30_5 ( );
FILL FILL_30_6 ( );
FILL FILL_30_7 ( );
FILL FILL_30_0_0 ( );
FILL FILL_30_0_1 ( );
FILL FILL_30_0_2 ( );
FILL FILL_30_1_0 ( );
FILL FILL_30_1_1 ( );
FILL FILL_30_1_2 ( );
FILL FILL_30_2_0 ( );
FILL FILL_30_2_1 ( );
FILL FILL_30_2_2 ( );
FILL FILL_30_3_0 ( );
FILL FILL_30_3_1 ( );
FILL FILL_30_3_2 ( );
FILL FILL_30_4_0 ( );
FILL FILL_30_4_1 ( );
FILL FILL_30_4_2 ( );
FILL FILL_30_5_0 ( );
FILL FILL_30_5_1 ( );
FILL FILL_30_5_2 ( );
FILL FILL_30_6_0 ( );
FILL FILL_30_6_1 ( );
FILL FILL_30_6_2 ( );
FILL FILL_31_1 ( );
FILL FILL_31_2 ( );
FILL FILL_31_3 ( );
FILL FILL_31_4 ( );
FILL FILL_31_5 ( );
FILL FILL_31_6 ( );
FILL FILL_31_0_0 ( );
FILL FILL_31_0_1 ( );
FILL FILL_31_0_2 ( );
FILL FILL_31_1_0 ( );
FILL FILL_31_1_1 ( );
FILL FILL_31_1_2 ( );
FILL FILL_31_2_0 ( );
FILL FILL_31_2_1 ( );
FILL FILL_31_2_2 ( );
FILL FILL_31_3_0 ( );
FILL FILL_31_3_1 ( );
FILL FILL_31_3_2 ( );
FILL FILL_31_4_0 ( );
FILL FILL_31_4_1 ( );
FILL FILL_31_4_2 ( );
FILL FILL_31_5_0 ( );
FILL FILL_31_5_1 ( );
FILL FILL_31_5_2 ( );
FILL FILL_31_6_0 ( );
FILL FILL_31_6_1 ( );
FILL FILL_31_6_2 ( );
FILL FILL_32_1 ( );
FILL FILL_32_2 ( );
FILL FILL_32_3 ( );
FILL FILL_32_0_0 ( );
FILL FILL_32_0_1 ( );
FILL FILL_32_0_2 ( );
FILL FILL_32_1_0 ( );
FILL FILL_32_1_1 ( );
FILL FILL_32_1_2 ( );
FILL FILL_32_2_0 ( );
FILL FILL_32_2_1 ( );
FILL FILL_32_2_2 ( );
FILL FILL_32_3_0 ( );
FILL FILL_32_3_1 ( );
FILL FILL_32_3_2 ( );
FILL FILL_32_4_0 ( );
FILL FILL_32_4_1 ( );
FILL FILL_32_4_2 ( );
FILL FILL_32_5_0 ( );
FILL FILL_32_5_1 ( );
FILL FILL_32_5_2 ( );
FILL FILL_32_6_0 ( );
FILL FILL_32_6_1 ( );
FILL FILL_32_6_2 ( );
FILL FILL_33_1 ( );
FILL FILL_33_2 ( );
FILL FILL_33_0_0 ( );
FILL FILL_33_0_1 ( );
FILL FILL_33_0_2 ( );
FILL FILL_33_1_0 ( );
FILL FILL_33_1_1 ( );
FILL FILL_33_1_2 ( );
FILL FILL_33_2_0 ( );
FILL FILL_33_2_1 ( );
FILL FILL_33_2_2 ( );
FILL FILL_33_3_0 ( );
FILL FILL_33_3_1 ( );
FILL FILL_33_3_2 ( );
FILL FILL_33_4_0 ( );
FILL FILL_33_4_1 ( );
FILL FILL_33_4_2 ( );
FILL FILL_33_5_0 ( );
FILL FILL_33_5_1 ( );
FILL FILL_33_5_2 ( );
FILL FILL_33_6_0 ( );
FILL FILL_33_6_1 ( );
FILL FILL_33_6_2 ( );
FILL FILL_34_1 ( );
FILL FILL_34_2 ( );
FILL FILL_34_3 ( );
FILL FILL_34_0_0 ( );
FILL FILL_34_0_1 ( );
FILL FILL_34_0_2 ( );
FILL FILL_34_1_0 ( );
FILL FILL_34_1_1 ( );
FILL FILL_34_1_2 ( );
FILL FILL_34_2_0 ( );
FILL FILL_34_2_1 ( );
FILL FILL_34_2_2 ( );
FILL FILL_34_3_0 ( );
FILL FILL_34_3_1 ( );
FILL FILL_34_3_2 ( );
FILL FILL_34_4_0 ( );
FILL FILL_34_4_1 ( );
FILL FILL_34_4_2 ( );
FILL FILL_34_5_0 ( );
FILL FILL_34_5_1 ( );
FILL FILL_34_5_2 ( );
FILL FILL_34_6_0 ( );
FILL FILL_34_6_1 ( );
FILL FILL_34_6_2 ( );
FILL FILL_35_1 ( );
FILL FILL_35_0_0 ( );
FILL FILL_35_0_1 ( );
FILL FILL_35_0_2 ( );
FILL FILL_35_1_0 ( );
FILL FILL_35_1_1 ( );
FILL FILL_35_1_2 ( );
FILL FILL_35_2_0 ( );
FILL FILL_35_2_1 ( );
FILL FILL_35_2_2 ( );
FILL FILL_35_3_0 ( );
FILL FILL_35_3_1 ( );
FILL FILL_35_3_2 ( );
FILL FILL_35_4_0 ( );
FILL FILL_35_4_1 ( );
FILL FILL_35_4_2 ( );
FILL FILL_35_5_0 ( );
FILL FILL_35_5_1 ( );
FILL FILL_35_5_2 ( );
FILL FILL_35_6_0 ( );
FILL FILL_35_6_1 ( );
FILL FILL_35_6_2 ( );
FILL FILL_36_1 ( );
FILL FILL_36_2 ( );
FILL FILL_36_3 ( );
FILL FILL_36_4 ( );
FILL FILL_36_5 ( );
FILL FILL_36_6 ( );
FILL FILL_36_0_0 ( );
FILL FILL_36_0_1 ( );
FILL FILL_36_0_2 ( );
FILL FILL_36_1_0 ( );
FILL FILL_36_1_1 ( );
FILL FILL_36_1_2 ( );
FILL FILL_36_2_0 ( );
FILL FILL_36_2_1 ( );
FILL FILL_36_2_2 ( );
FILL FILL_36_3_0 ( );
FILL FILL_36_3_1 ( );
FILL FILL_36_3_2 ( );
FILL FILL_36_4_0 ( );
FILL FILL_36_4_1 ( );
FILL FILL_36_4_2 ( );
FILL FILL_36_5_0 ( );
FILL FILL_36_5_1 ( );
FILL FILL_36_5_2 ( );
FILL FILL_36_6_0 ( );
FILL FILL_36_6_1 ( );
FILL FILL_36_6_2 ( );
FILL FILL_37_1 ( );
FILL FILL_37_2 ( );
FILL FILL_37_3 ( );
FILL FILL_37_4 ( );
FILL FILL_37_5 ( );
FILL FILL_37_0_0 ( );
FILL FILL_37_0_1 ( );
FILL FILL_37_0_2 ( );
FILL FILL_37_1_0 ( );
FILL FILL_37_1_1 ( );
FILL FILL_37_1_2 ( );
FILL FILL_37_2_0 ( );
FILL FILL_37_2_1 ( );
FILL FILL_37_2_2 ( );
FILL FILL_37_3_0 ( );
FILL FILL_37_3_1 ( );
FILL FILL_37_3_2 ( );
FILL FILL_37_4_0 ( );
FILL FILL_37_4_1 ( );
FILL FILL_37_4_2 ( );
FILL FILL_37_5_0 ( );
FILL FILL_37_5_1 ( );
FILL FILL_37_5_2 ( );
FILL FILL_37_6_0 ( );
FILL FILL_37_6_1 ( );
FILL FILL_37_6_2 ( );
FILL FILL_38_0_0 ( );
FILL FILL_38_0_1 ( );
FILL FILL_38_0_2 ( );
FILL FILL_38_1_0 ( );
FILL FILL_38_1_1 ( );
FILL FILL_38_1_2 ( );
FILL FILL_38_2_0 ( );
FILL FILL_38_2_1 ( );
FILL FILL_38_2_2 ( );
FILL FILL_38_3_0 ( );
FILL FILL_38_3_1 ( );
FILL FILL_38_3_2 ( );
FILL FILL_38_4_0 ( );
FILL FILL_38_4_1 ( );
FILL FILL_38_4_2 ( );
FILL FILL_38_5_0 ( );
FILL FILL_38_5_1 ( );
FILL FILL_38_5_2 ( );
FILL FILL_38_6_0 ( );
FILL FILL_38_6_1 ( );
FILL FILL_38_6_2 ( );
FILL FILL_39_1 ( );
FILL FILL_39_2 ( );
FILL FILL_39_3 ( );
FILL FILL_39_4 ( );
FILL FILL_39_0_0 ( );
FILL FILL_39_0_1 ( );
FILL FILL_39_0_2 ( );
FILL FILL_39_1_0 ( );
FILL FILL_39_1_1 ( );
FILL FILL_39_1_2 ( );
FILL FILL_39_2_0 ( );
FILL FILL_39_2_1 ( );
FILL FILL_39_2_2 ( );
FILL FILL_39_3_0 ( );
FILL FILL_39_3_1 ( );
FILL FILL_39_3_2 ( );
FILL FILL_39_4_0 ( );
FILL FILL_39_4_1 ( );
FILL FILL_39_4_2 ( );
FILL FILL_39_5_0 ( );
FILL FILL_39_5_1 ( );
FILL FILL_39_5_2 ( );
FILL FILL_39_6_0 ( );
FILL FILL_39_6_1 ( );
FILL FILL_39_6_2 ( );
FILL FILL_40_0_0 ( );
FILL FILL_40_0_1 ( );
FILL FILL_40_0_2 ( );
FILL FILL_40_1_0 ( );
FILL FILL_40_1_1 ( );
FILL FILL_40_1_2 ( );
FILL FILL_40_2_0 ( );
FILL FILL_40_2_1 ( );
FILL FILL_40_2_2 ( );
FILL FILL_40_3_0 ( );
FILL FILL_40_3_1 ( );
FILL FILL_40_3_2 ( );
FILL FILL_40_4_0 ( );
FILL FILL_40_4_1 ( );
FILL FILL_40_4_2 ( );
FILL FILL_40_5_0 ( );
FILL FILL_40_5_1 ( );
FILL FILL_40_5_2 ( );
FILL FILL_40_6_0 ( );
FILL FILL_40_6_1 ( );
FILL FILL_40_6_2 ( );
FILL FILL_41_0_0 ( );
FILL FILL_41_0_1 ( );
FILL FILL_41_0_2 ( );
FILL FILL_41_1_0 ( );
FILL FILL_41_1_1 ( );
FILL FILL_41_1_2 ( );
FILL FILL_41_2_0 ( );
FILL FILL_41_2_1 ( );
FILL FILL_41_2_2 ( );
FILL FILL_41_3_0 ( );
FILL FILL_41_3_1 ( );
FILL FILL_41_3_2 ( );
FILL FILL_41_4_0 ( );
FILL FILL_41_4_1 ( );
FILL FILL_41_4_2 ( );
FILL FILL_41_5_0 ( );
FILL FILL_41_5_1 ( );
FILL FILL_41_5_2 ( );
FILL FILL_41_6_0 ( );
FILL FILL_41_6_1 ( );
FILL FILL_41_6_2 ( );
FILL FILL_42_1 ( );
FILL FILL_42_2 ( );
FILL FILL_42_3 ( );
FILL FILL_42_4 ( );
FILL FILL_42_5 ( );
FILL FILL_42_0_0 ( );
FILL FILL_42_0_1 ( );
FILL FILL_42_0_2 ( );
FILL FILL_42_1_0 ( );
FILL FILL_42_1_1 ( );
FILL FILL_42_1_2 ( );
FILL FILL_42_2_0 ( );
FILL FILL_42_2_1 ( );
FILL FILL_42_2_2 ( );
FILL FILL_42_3_0 ( );
FILL FILL_42_3_1 ( );
FILL FILL_42_3_2 ( );
FILL FILL_42_4_0 ( );
FILL FILL_42_4_1 ( );
FILL FILL_42_4_2 ( );
FILL FILL_42_5_0 ( );
FILL FILL_42_5_1 ( );
FILL FILL_42_5_2 ( );
FILL FILL_42_6_0 ( );
FILL FILL_42_6_1 ( );
FILL FILL_42_6_2 ( );
FILL FILL_43_1 ( );
FILL FILL_43_0_0 ( );
FILL FILL_43_0_1 ( );
FILL FILL_43_0_2 ( );
FILL FILL_43_1_0 ( );
FILL FILL_43_1_1 ( );
FILL FILL_43_1_2 ( );
FILL FILL_43_2_0 ( );
FILL FILL_43_2_1 ( );
FILL FILL_43_2_2 ( );
FILL FILL_43_3_0 ( );
FILL FILL_43_3_1 ( );
FILL FILL_43_3_2 ( );
FILL FILL_43_4_0 ( );
FILL FILL_43_4_1 ( );
FILL FILL_43_4_2 ( );
FILL FILL_43_5_0 ( );
FILL FILL_43_5_1 ( );
FILL FILL_43_5_2 ( );
FILL FILL_43_6_0 ( );
FILL FILL_43_6_1 ( );
FILL FILL_43_6_2 ( );
FILL FILL_44_1 ( );
FILL FILL_44_2 ( );
FILL FILL_44_3 ( );
FILL FILL_44_4 ( );
FILL FILL_44_5 ( );
FILL FILL_44_6 ( );
FILL FILL_44_0_0 ( );
FILL FILL_44_0_1 ( );
FILL FILL_44_0_2 ( );
FILL FILL_44_1_0 ( );
FILL FILL_44_1_1 ( );
FILL FILL_44_1_2 ( );
FILL FILL_44_2_0 ( );
FILL FILL_44_2_1 ( );
FILL FILL_44_2_2 ( );
FILL FILL_44_3_0 ( );
FILL FILL_44_3_1 ( );
FILL FILL_44_3_2 ( );
FILL FILL_44_4_0 ( );
FILL FILL_44_4_1 ( );
FILL FILL_44_4_2 ( );
FILL FILL_44_5_0 ( );
FILL FILL_44_5_1 ( );
FILL FILL_44_5_2 ( );
FILL FILL_44_6_0 ( );
FILL FILL_44_6_1 ( );
FILL FILL_44_6_2 ( );
FILL FILL_45_1 ( );
FILL FILL_45_2 ( );
FILL FILL_45_0_0 ( );
FILL FILL_45_0_1 ( );
FILL FILL_45_0_2 ( );
FILL FILL_45_1_0 ( );
FILL FILL_45_1_1 ( );
FILL FILL_45_1_2 ( );
FILL FILL_45_2_0 ( );
FILL FILL_45_2_1 ( );
FILL FILL_45_2_2 ( );
FILL FILL_45_3_0 ( );
FILL FILL_45_3_1 ( );
FILL FILL_45_3_2 ( );
FILL FILL_45_4_0 ( );
FILL FILL_45_4_1 ( );
FILL FILL_45_4_2 ( );
FILL FILL_45_5_0 ( );
FILL FILL_45_5_1 ( );
FILL FILL_45_5_2 ( );
FILL FILL_45_6_0 ( );
FILL FILL_45_6_1 ( );
FILL FILL_45_6_2 ( );
FILL FILL_46_1 ( );
FILL FILL_46_2 ( );
FILL FILL_46_3 ( );
FILL FILL_46_0_0 ( );
FILL FILL_46_0_1 ( );
FILL FILL_46_0_2 ( );
FILL FILL_46_1_0 ( );
FILL FILL_46_1_1 ( );
FILL FILL_46_1_2 ( );
FILL FILL_46_2_0 ( );
FILL FILL_46_2_1 ( );
FILL FILL_46_2_2 ( );
FILL FILL_46_3_0 ( );
FILL FILL_46_3_1 ( );
FILL FILL_46_3_2 ( );
FILL FILL_46_4_0 ( );
FILL FILL_46_4_1 ( );
FILL FILL_46_4_2 ( );
FILL FILL_46_5_0 ( );
FILL FILL_46_5_1 ( );
FILL FILL_46_5_2 ( );
FILL FILL_46_6_0 ( );
FILL FILL_46_6_1 ( );
FILL FILL_46_6_2 ( );
FILL FILL_47_1 ( );
FILL FILL_47_2 ( );
FILL FILL_47_3 ( );
FILL FILL_47_0_0 ( );
FILL FILL_47_0_1 ( );
FILL FILL_47_0_2 ( );
FILL FILL_47_1_0 ( );
FILL FILL_47_1_1 ( );
FILL FILL_47_1_2 ( );
FILL FILL_47_2_0 ( );
FILL FILL_47_2_1 ( );
FILL FILL_47_2_2 ( );
FILL FILL_47_3_0 ( );
FILL FILL_47_3_1 ( );
FILL FILL_47_3_2 ( );
FILL FILL_47_4_0 ( );
FILL FILL_47_4_1 ( );
FILL FILL_47_4_2 ( );
FILL FILL_47_5_0 ( );
FILL FILL_47_5_1 ( );
FILL FILL_47_5_2 ( );
FILL FILL_47_6_0 ( );
FILL FILL_47_6_1 ( );
FILL FILL_47_6_2 ( );
FILL FILL_48_1 ( );
FILL FILL_48_2 ( );
FILL FILL_48_3 ( );
FILL FILL_48_4 ( );
FILL FILL_48_5 ( );
FILL FILL_48_6 ( );
FILL FILL_48_0_0 ( );
FILL FILL_48_0_1 ( );
FILL FILL_48_0_2 ( );
FILL FILL_48_1_0 ( );
FILL FILL_48_1_1 ( );
FILL FILL_48_1_2 ( );
FILL FILL_48_2_0 ( );
FILL FILL_48_2_1 ( );
FILL FILL_48_2_2 ( );
FILL FILL_48_3_0 ( );
FILL FILL_48_3_1 ( );
FILL FILL_48_3_2 ( );
FILL FILL_48_4_0 ( );
FILL FILL_48_4_1 ( );
FILL FILL_48_4_2 ( );
FILL FILL_48_5_0 ( );
FILL FILL_48_5_1 ( );
FILL FILL_48_5_2 ( );
FILL FILL_48_6_0 ( );
FILL FILL_48_6_1 ( );
FILL FILL_48_6_2 ( );
FILL FILL_49_1 ( );
FILL FILL_49_2 ( );
FILL FILL_49_3 ( );
FILL FILL_49_4 ( );
FILL FILL_49_5 ( );
FILL FILL_49_6 ( );
FILL FILL_49_7 ( );
FILL FILL_49_8 ( );
FILL FILL_49_9 ( );
FILL FILL_49_0_0 ( );
FILL FILL_49_0_1 ( );
FILL FILL_49_0_2 ( );
FILL FILL_49_1_0 ( );
FILL FILL_49_1_1 ( );
FILL FILL_49_1_2 ( );
FILL FILL_49_2_0 ( );
FILL FILL_49_2_1 ( );
FILL FILL_49_2_2 ( );
FILL FILL_49_3_0 ( );
FILL FILL_49_3_1 ( );
FILL FILL_49_3_2 ( );
FILL FILL_49_4_0 ( );
FILL FILL_49_4_1 ( );
FILL FILL_49_4_2 ( );
FILL FILL_49_5_0 ( );
FILL FILL_49_5_1 ( );
FILL FILL_49_5_2 ( );
FILL FILL_49_6_0 ( );
FILL FILL_49_6_1 ( );
FILL FILL_49_6_2 ( );
FILL FILL_50_1 ( );
FILL FILL_50_2 ( );
FILL FILL_50_3 ( );
FILL FILL_50_4 ( );
FILL FILL_50_5 ( );
FILL FILL_50_6 ( );
FILL FILL_50_7 ( );
FILL FILL_50_8 ( );
FILL FILL_50_9 ( );
FILL FILL_50_0_0 ( );
FILL FILL_50_0_1 ( );
FILL FILL_50_0_2 ( );
FILL FILL_50_1_0 ( );
FILL FILL_50_1_1 ( );
FILL FILL_50_1_2 ( );
FILL FILL_50_2_0 ( );
FILL FILL_50_2_1 ( );
FILL FILL_50_2_2 ( );
FILL FILL_50_3_0 ( );
FILL FILL_50_3_1 ( );
FILL FILL_50_3_2 ( );
FILL FILL_50_4_0 ( );
FILL FILL_50_4_1 ( );
FILL FILL_50_4_2 ( );
FILL FILL_50_5_0 ( );
FILL FILL_50_5_1 ( );
FILL FILL_50_5_2 ( );
FILL FILL_50_6_0 ( );
FILL FILL_50_6_1 ( );
FILL FILL_50_6_2 ( );
FILL FILL_51_1 ( );
FILL FILL_51_2 ( );
FILL FILL_51_3 ( );
FILL FILL_51_4 ( );
FILL FILL_51_5 ( );
FILL FILL_51_0_0 ( );
FILL FILL_51_0_1 ( );
FILL FILL_51_0_2 ( );
FILL FILL_51_1_0 ( );
FILL FILL_51_1_1 ( );
FILL FILL_51_1_2 ( );
FILL FILL_51_2_0 ( );
FILL FILL_51_2_1 ( );
FILL FILL_51_2_2 ( );
FILL FILL_51_3_0 ( );
FILL FILL_51_3_1 ( );
FILL FILL_51_3_2 ( );
FILL FILL_51_4_0 ( );
FILL FILL_51_4_1 ( );
FILL FILL_51_4_2 ( );
FILL FILL_51_5_0 ( );
FILL FILL_51_5_1 ( );
FILL FILL_51_5_2 ( );
FILL FILL_51_6_0 ( );
FILL FILL_51_6_1 ( );
FILL FILL_51_6_2 ( );
FILL FILL_52_1 ( );
FILL FILL_52_2 ( );
FILL FILL_52_0_0 ( );
FILL FILL_52_0_1 ( );
FILL FILL_52_0_2 ( );
FILL FILL_52_1_0 ( );
FILL FILL_52_1_1 ( );
FILL FILL_52_1_2 ( );
FILL FILL_52_2_0 ( );
FILL FILL_52_2_1 ( );
FILL FILL_52_2_2 ( );
FILL FILL_52_3_0 ( );
FILL FILL_52_3_1 ( );
FILL FILL_52_3_2 ( );
FILL FILL_52_4_0 ( );
FILL FILL_52_4_1 ( );
FILL FILL_52_4_2 ( );
FILL FILL_52_5_0 ( );
FILL FILL_52_5_1 ( );
FILL FILL_52_5_2 ( );
FILL FILL_52_6_0 ( );
FILL FILL_52_6_1 ( );
FILL FILL_52_6_2 ( );
FILL FILL_53_1 ( );
FILL FILL_53_2 ( );
FILL FILL_53_3 ( );
FILL FILL_53_4 ( );
FILL FILL_53_5 ( );
FILL FILL_53_0_0 ( );
FILL FILL_53_0_1 ( );
FILL FILL_53_0_2 ( );
FILL FILL_53_1_0 ( );
FILL FILL_53_1_1 ( );
FILL FILL_53_1_2 ( );
FILL FILL_53_2_0 ( );
FILL FILL_53_2_1 ( );
FILL FILL_53_2_2 ( );
FILL FILL_53_3_0 ( );
FILL FILL_53_3_1 ( );
FILL FILL_53_3_2 ( );
FILL FILL_53_4_0 ( );
FILL FILL_53_4_1 ( );
FILL FILL_53_4_2 ( );
FILL FILL_53_5_0 ( );
FILL FILL_53_5_1 ( );
FILL FILL_53_5_2 ( );
FILL FILL_53_6_0 ( );
FILL FILL_53_6_1 ( );
FILL FILL_53_6_2 ( );
FILL FILL_54_1 ( );
FILL FILL_54_2 ( );
FILL FILL_54_3 ( );
FILL FILL_54_4 ( );
FILL FILL_54_5 ( );
FILL FILL_54_6 ( );
FILL FILL_54_7 ( );
FILL FILL_54_8 ( );
FILL FILL_54_0_0 ( );
FILL FILL_54_0_1 ( );
FILL FILL_54_0_2 ( );
FILL FILL_54_1_0 ( );
FILL FILL_54_1_1 ( );
FILL FILL_54_1_2 ( );
FILL FILL_54_2_0 ( );
FILL FILL_54_2_1 ( );
FILL FILL_54_2_2 ( );
FILL FILL_54_3_0 ( );
FILL FILL_54_3_1 ( );
FILL FILL_54_3_2 ( );
FILL FILL_54_4_0 ( );
FILL FILL_54_4_1 ( );
FILL FILL_54_4_2 ( );
FILL FILL_54_5_0 ( );
FILL FILL_54_5_1 ( );
FILL FILL_54_5_2 ( );
FILL FILL_54_6_0 ( );
FILL FILL_54_6_1 ( );
FILL FILL_54_6_2 ( );
FILL FILL_55_1 ( );
FILL FILL_55_2 ( );
FILL FILL_55_3 ( );
FILL FILL_55_4 ( );
FILL FILL_55_5 ( );
FILL FILL_55_6 ( );
FILL FILL_55_7 ( );
FILL FILL_55_8 ( );
FILL FILL_55_9 ( );
FILL FILL_55_10 ( );
endmodule

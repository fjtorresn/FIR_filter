* NGSPICE file created from fir2n.ext - technology: scmos

* Black-box entry subcircuit for FILL abstract view
.subckt FILL gnd vdd
.ends

* Black-box entry subcircuit for NAND3X1 abstract view
.subckt NAND3X1 A B C gnd Y vdd
.ends

* Black-box entry subcircuit for NOR2X1 abstract view
.subckt NOR2X1 A B gnd Y vdd
.ends

* Black-box entry subcircuit for CLKBUF1 abstract view
.subckt CLKBUF1 A gnd Y vdd
.ends

* Black-box entry subcircuit for OAI21X1 abstract view
.subckt OAI21X1 A B C gnd Y vdd
.ends

* Black-box entry subcircuit for BUFX2 abstract view
.subckt BUFX2 A gnd Y vdd
.ends

* Black-box entry subcircuit for NAND2X1 abstract view
.subckt NAND2X1 A B gnd Y vdd
.ends

* Black-box entry subcircuit for AOI21X1 abstract view
.subckt AOI21X1 A B C gnd Y vdd
.ends

* Black-box entry subcircuit for DFFPOSX1 abstract view
.subckt DFFPOSX1 Q CLK D gnd vdd
.ends

* Black-box entry subcircuit for DFFSR abstract view
.subckt DFFSR Q CLK R S D gnd vdd
.ends

* Black-box entry subcircuit for AOI22X1 abstract view
.subckt AOI22X1 A B C D gnd Y vdd
.ends

* Black-box entry subcircuit for OAI22X1 abstract view
.subckt OAI22X1 A B C D gnd Y vdd
.ends

* Black-box entry subcircuit for INVX1 abstract view
.subckt INVX1 A gnd Y vdd
.ends

* Black-box entry subcircuit for AND2X2 abstract view
.subckt AND2X2 A B gnd Y vdd
.ends

* Black-box entry subcircuit for XOR2X1 abstract view
.subckt XOR2X1 A B gnd Y vdd
.ends

* Black-box entry subcircuit for OR2X2 abstract view
.subckt OR2X2 A B gnd Y vdd
.ends

* Black-box entry subcircuit for NOR3X1 abstract view
.subckt NOR3X1 A B C gnd Y vdd
.ends

* Black-box entry subcircuit for XNOR2X1 abstract view
.subckt XNOR2X1 A B gnd Y vdd
.ends

.subckt fir2n clk rst din[0] din[1] din[2] din[3] din[4] din[5] din[6] din[7] dout[0]
+ dout[1] dout[2] dout[3] dout[4] dout[5] dout[6] dout[7]
XFILL_22_DFFSR_143 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_8_CLKBUF1_8 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_2_DFFSR_25 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_36_DFFSR_247 BUFX2_99/A DFFSR_7/S FILL
XFILL_19_DFFSR_18 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_12_DFFSR_146 BUFX2_79/A DFFSR_7/S FILL
XFILL_6_BUFX2_53 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_26_DFFSR_250 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_16_DFFSR_253 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_1_NOR2X1_6 BUFX2_98/A DFFSR_6/S FILL
XFILL_6_NAND3X1_172 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_19_CLKBUF1_11 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_43_DFFSR_75 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_8_DFFSR_140 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_40_2_0 BUFX2_98/A DFFSR_6/S FILL
XFILL_49_DFFSR_171 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_18_CLKBUF1_14 DFFSR_34/gnd DFFSR_34/S FILL
XNAND3X1_208 NAND3X1_214/A NAND3X1_214/B OAI21X1_59/Y DFFSR_46/gnd XOR2X1_8/A DFFSR_54/S
+ NAND3X1
XFILL_1_INVX1_117 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_39_DFFSR_174 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_17_CLKBUF1_17 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_27_DFFSR_25 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_16_DFFSR_65 BUFX2_79/A DFFSR_7/S FILL
XFILL_38_4_1 BUFX2_79/A DFFSR_7/S FILL
XFILL_7_NAND3X1_106 INVX1_3/gnd DFFSR_23/S FILL
XFILL_2_DFFSR_250 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_16_CLKBUF1_20 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_29_DFFSR_177 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_11_DFFPOSX1_10 INVX1_67/gnd DFFSR_201/S FILL
XFILL_15_CLKBUF1_23 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_19_DFFSR_180 DFFSR_34/gnd DFFSR_34/S FILL
XNOR2X1_62 BUFX2_7/Y BUFX2_36/Y INVX1_67/gnd NOR2X1_62/Y DFFSR_201/S NOR2X1
XFILL_36_6_2 BUFX2_99/A DFFSR_92/S FILL
XFILL_14_CLKBUF1_26 INVX1_1/gnd DFFSR_53/S FILL
XFILL_3_XOR2X1_2 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_23_DFFSR_4 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_13_CLKBUF1_29 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_4_NOR2X1_59 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_6_OAI21X1_7 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_12_CLKBUF1_32 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_42_DFFSR_101 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_35_DFFSR_32 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_7_DFFSR_79 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_24_DFFSR_72 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_11_CLKBUF1_35 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_5_DFFSR_177 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_32_DFFSR_104 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_10_CLKBUF1_38 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_5_NAND3X1_202 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_46_DFFSR_208 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_22_DFFSR_107 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_36_DFFSR_211 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_1_DFFPOSX1_21 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_1_AND2X2_21 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_12_DFFSR_110 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_6_BUFX2_17 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_26_DFFSR_214 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_9_CLKBUF1_41 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_16_DFFSR_217 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_8_CLKBUF1_44 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_6_NAND3X1_136 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_7_CLKBUF1_47 BUFX2_98/A DFFSR_32/S FILL
XFILL_10_DFFPOSX1_40 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_8_DFFSR_104 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_32_DFFSR_79 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_43_DFFSR_39 INVX1_3/gnd DFFSR_79/S FILL
XFILL_4_INVX1_73 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_49_DFFSR_135 DFFSR_62/gnd DFFSR_208/S FILL
XNAND3X1_172 INVX1_158/A OAI21X1_48/Y OAI21X1_49/Y DFFSR_1/gnd AOI22X1_23/B DFFSR_1/S
+ NAND3X1
XFILL_39_DFFSR_138 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_16_DFFSR_29 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_2_DFFSR_214 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_3_BUFX2_64 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_29_DFFSR_141 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_46_1_2 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_43_DFFSR_245 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_20_DFFPOSX1_29 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_5_CLKBUF1_9 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_19_DFFSR_144 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_33_DFFSR_248 DFFSR_28/gnd DFFSR_8/S FILL
XNOR2X1_26 NOR2X1_26/A NOR2X1_26/B DFFSR_8/gnd NOR2X1_26/Y DFFSR_60/S NOR2X1
XFILL_23_DFFSR_251 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_4_NAND3X1_232 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_40_DFFSR_86 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_4_NOR2X1_23 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_13_DFFSR_254 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_7_DFFSR_43 BUFX2_98/A DFFSR_6/S FILL
XFILL_24_DFFSR_36 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_13_DFFSR_76 BUFX2_79/A DFFSR_7/S FILL
XFILL_5_DFFSR_141 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_5_NAND3X1_166 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_14_0_0 INVX1_39/gnd DFFSR_54/S FILL
XFILL_46_DFFSR_172 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_9_DFFSR_248 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_36_DFFSR_175 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_50_DFFSR_279 BUFX2_99/A DFFSR_7/S FILL
XFILL_26_DFFSR_178 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_12_2_1 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_48_DFFSR_93 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_16_DFFSR_181 INVX1_3/gnd DFFSR_79/S FILL
XFILL_6_NAND3X1_100 AND2X2_38/B DFFSR_59/S FILL
XFILL_7_CLKBUF1_11 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_9_AND2X2_2 BUFX2_99/A DFFSR_7/S FILL
XFILL_10_4_2 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_4_DFFSR_90 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_4_INVX1_37 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_32_DFFSR_43 BUFX2_98/A DFFSR_6/S FILL
XFILL_21_DFFSR_83 INVX1_3/gnd DFFSR_79/S FILL
XFILL_1_NOR2X1_60 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_6_CLKBUF1_14 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_3_OAI21X1_8 BUFX2_99/A DFFSR_7/S FILL
XFILL_5_CLKBUF1_17 BUFX2_8/gnd DFFSR_81/S FILL
XNAND3X1_136 NOR3X1_1/A INVX1_130/Y AND2X2_28/Y DFFSR_1/gnd AOI21X1_6/A DFFSR_81/S
+ NAND3X1
XFILL_39_DFFSR_102 DFFSR_4/gnd DFFSR_98/S FILL
XCLKBUF1_14 BUFX2_5/Y DFFSR_34/gnd CLKBUF1_14/Y DFFSR_34/S CLKBUF1
XFILL_5_4 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_4_CLKBUF1_20 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_2_DFFSR_178 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_3_BUFX2_28 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_29_DFFSR_105 INVX1_1/gnd DFFSR_53/S FILL
XFILL_43_DFFSR_209 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_3_CLKBUF1_23 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_8_AND2X2_19 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_19_DFFSR_108 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_6_OAI21X1_118 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_33_DFFSR_212 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_2_CLKBUF1_26 INVX1_1/gnd DFFSR_53/S FILL
XFILL_23_DFFSR_215 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_1_CLKBUF1_29 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_4_NAND3X1_196 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_40_DFFSR_50 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_1_INVX1_84 INVX1_39/gnd DFFSR_34/S FILL
XFILL_29_DFFSR_90 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_0_DFFPOSX1_15 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_13_DFFSR_218 BUFX2_98/A DFFSR_32/S FILL
XFILL_0_CLKBUF1_32 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_13_DFFSR_40 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_5_DFFSR_105 INVX1_1/gnd DFFSR_53/S FILL
XFILL_0_BUFX2_75 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_46_DFFSR_136 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_5_NAND3X1_130 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_9_DFFSR_212 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_36_DFFSR_139 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_50_DFFSR_243 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_26_DFFSR_142 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_35_DFFSR_7 BUFX2_79/A DFFSR_7/S FILL
XFILL_2_INVX1_189 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_40_DFFSR_246 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_48_DFFSR_57 BUFX2_79/A DFFSR_6/S FILL
XFILL_37_DFFSR_97 INVX1_1/gnd DFFSR_97/S FILL
XFILL_16_DFFSR_145 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_30_DFFSR_249 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_20_DFFSR_252 AND2X2_38/B DFFSR_23/S FILL
XFILL_21_DFFSR_47 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_19_DFFPOSX1_23 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_4_DFFSR_54 INVX1_39/gnd DFFSR_54/S FILL
XFILL_1_NOR2X1_24 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_10_DFFSR_87 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_10_DFFSR_255 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_0_0_2 BUFX2_72/gnd DFFSR_276/S FILL
XNAND3X1_100 NAND2X1_46/Y NAND3X1_97/Y AND2X2_23/Y AND2X2_38/B NOR2X1_49/A DFFSR_59/S
+ NAND3X1
XFILL_3_NAND3X1_226 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_2_DFFSR_142 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_43_DFFSR_173 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_6_DFFSR_249 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_33_DFFSR_176 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_47_DFFSR_280 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_23_DFFSR_179 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_4_NAND3X1_160 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_1_INVX1_48 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_40_DFFSR_14 INVX1_1/gnd DFFSR_53/S FILL
XFILL_18_DFFSR_94 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_29_DFFSR_54 INVX1_39/gnd DFFSR_54/S FILL
XFILL_13_DFFSR_182 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_47_2_0 DFFSR_8/gnd DFFSR_60/S FILL
XOAI21X1_118 XOR2X1_15/Y OR2X2_6/Y INVX1_212/Y OR2X2_6/gnd AOI21X1_70/C DFFSR_53/S
+ OAI21X1
XFILL_9_DFFPOSX1_34 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_0_BUFX2_39 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_45_4_1 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_0_OAI21X1_9 INVX1_67/gnd DFFSR_201/S FILL
XFILL_46_DFFSR_100 INVX1_1/gnd DFFSR_97/S FILL
XFILL_9_DFFSR_176 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_36_DFFSR_103 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_50_DFFSR_207 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_43_6_2 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_26_DFFSR_106 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_2_INVX1_153 INVX1_67/gnd DFFSR_175/S FILL
XFILL_40_DFFSR_210 BUFX2_98/A DFFSR_6/S FILL
XFILL_37_DFFSR_61 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_48_DFFSR_21 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_5_AND2X2_20 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_16_DFFSR_109 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_30_DFFSR_213 INVX1_3/gnd DFFSR_23/S FILL
XFILL_20_DFFSR_216 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_4_DFFSR_18 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_21_DFFSR_11 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_10_DFFSR_51 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_5_OAI21X1_112 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_10_DFFSR_219 INVX1_67/gnd DFFSR_175/S FILL
XFILL_3_NAND3X1_190 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_2_DFFSR_106 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_11_5_0 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_43_DFFSR_137 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_22_DFFSR_1 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_45_DFFSR_68 BUFX2_98/A DFFSR_6/S FILL
XFILL_6_DFFSR_213 INVX1_3/gnd DFFSR_23/S FILL
XFILL_33_DFFSR_140 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_47_DFFSR_244 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_23_DFFSR_143 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_9_CLKBUF1_8 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_4_NAND3X1_124 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_1_INVX1_12 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_1_DFFSR_65 BUFX2_79/A DFFSR_7/S FILL
XFILL_37_DFFSR_247 BUFX2_99/A DFFSR_7/S FILL
XFILL_18_DFFSR_58 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_29_DFFSR_18 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_13_DFFSR_146 BUFX2_79/A DFFSR_7/S FILL
XFILL_5_BUFX2_93 AND2X2_38/B DFFSR_59/S FILL
XFILL_27_DFFSR_250 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_6_BUFX2_2 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_6_NAND2X1_160 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_49_5 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_17_DFFSR_253 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_53_1_2 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_9_DFFSR_140 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_18_DFFPOSX1_17 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_50_DFFSR_171 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_2_INVX1_117 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_40_DFFSR_174 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_9_DFFSR_72 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_37_DFFSR_25 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_26_DFFSR_65 BUFX2_79/A DFFSR_7/S FILL
XFILL_2_NAND3X1_220 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_3_DFFSR_250 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_18_DFFPOSX1_2 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_30_DFFSR_177 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_17_DFFPOSX1_5 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_20_DFFSR_180 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_10_DFFSR_15 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_16_DFFPOSX1_8 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_10_DFFSR_183 INVX1_67/gnd DFFSR_175/S FILL
XFILL_3_NAND3X1_154 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_21_0_0 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_5_NOR2X1_59 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_7_OAI21X1_7 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_8_DFFPOSX1_28 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_43_DFFSR_101 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_45_DFFSR_32 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_34_DFFSR_72 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_19_2_1 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_6_DFFSR_177 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_33_DFFSR_104 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_47_DFFSR_208 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_1_1_0 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_23_DFFSR_107 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_37_DFFSR_211 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_1_DFFSR_29 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_18_DFFSR_22 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_17_4_2 DFFSR_34/gnd DFFSR_1/S FILL
XBUFX2_97 BUFX2_97/A OR2X2_3/gnd BUFX2_97/Y DFFSR_60/S BUFX2
XFILL_2_AND2X2_21 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_13_DFFSR_110 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_5_BUFX2_57 AND2X2_38/B DFFSR_23/S FILL
XFILL_27_DFFSR_214 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_17_DFFPOSX1_47 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_10_OAI22X1_3 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_6_NAND2X1_124 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_17_DFFSR_217 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_9_NOR3X1_3 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_9_DFFSR_104 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_42_DFFSR_79 NOR3X1_6/gnd DFFSR_79/S FILL
XNAND2X1_160 NAND2X1_160/A INVX1_208/Y NOR3X1_6/gnd AOI21X1_56/A DFFSR_79/S NAND2X1
XFILL_50_DFFSR_135 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_4_OAI21X1_106 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_27_DFFPOSX1_36 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_8_AOI21X1_52 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_40_DFFSR_138 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_26_DFFSR_29 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_9_DFFSR_36 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_7_AOI21X1_55 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_15_DFFSR_69 BUFX2_98/A DFFSR_32/S FILL
XFILL_2_NAND3X1_184 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_3_DFFSR_214 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_30_DFFSR_141 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_6_AOI21X1_58 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_44_DFFSR_245 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_6_CLKBUF1_9 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_20_DFFSR_144 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_34_DFFSR_248 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_5_AOI21X1_61 AND2X2_38/B DFFSR_59/S FILL
XAOI21X1_58 AOI21X1_58/A AOI21X1_58/B BUFX2_36/Y OR2X2_2/gnd AOI21X1_58/Y DFFSR_175/S
+ AOI21X1
XFILL_10_DFFSR_147 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_2_XOR2X1_6 BUFX2_99/A DFFSR_7/S FILL
XFILL_4_AOI21X1_64 AND2X2_38/B DFFSR_59/S FILL
XFILL_24_DFFSR_251 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_5_NOR2X1_23 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_13_DFFSR_8 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_50_DFFSR_86 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_3_NAND3X1_118 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_3_AOI21X1_67 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_14_DFFSR_254 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_2_AOI21X1_70 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_5_NAND2X1_154 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_6_DFFSR_83 INVX1_3/gnd DFFSR_79/S FILL
XFILL_34_DFFSR_36 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_23_DFFSR_76 BUFX2_79/A DFFSR_7/S FILL
XFILL_6_DFFSR_141 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_47_DFFSR_172 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_37_DFFSR_175 OR2X2_2/gnd DFFSR_175/S FILL
XBUFX2_61 BUFX2_60/A AND2X2_38/B BUFX2_61/Y DFFSR_59/S BUFX2
XFILL_0_DFFSR_251 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_5_BUFX2_21 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_17_DFFPOSX1_11 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_27_DFFSR_178 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_9_OAI21X1_97 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_7_0_2 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_17_DFFSR_181 INVX1_3/gnd DFFSR_79/S FILL
XFILL_34_DFFSR_4 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_1_NAND3X1_214 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_42_DFFSR_43 BUFX2_98/A DFFSR_6/S FILL
XFILL_31_DFFSR_83 INVX1_3/gnd DFFSR_79/S FILL
XFILL_3_INVX1_77 DFFSR_1/gnd DFFSR_81/S FILL
XNAND2X1_124 NAND2X1_59/A BUFX2_54/Y OR2X2_2/gnd OAI21X1_93/C DFFSR_216/S NAND2X1
XFILL_2_NOR2X1_60 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_4_OAI21X1_8 BUFX2_99/A DFFSR_7/S FILL
XFILL_8_AOI21X1_16 INVX1_67/gnd DFFSR_175/S FILL
XFILL_40_DFFSR_102 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_9_1 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_6_DFFPOSX1_2 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_7_AOI21X1_19 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_15_DFFSR_33 BUFX2_98/A DFFSR_32/S FILL
XFILL_2_NAND3X1_148 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_3_DFFSR_178 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_30_DFFSR_105 INVX1_1/gnd DFFSR_53/S FILL
XFILL_2_BUFX2_68 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_5_DFFPOSX1_5 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_6_AOI21X1_22 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_44_DFFSR_209 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_9_AND2X2_19 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_54_2_0 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_20_DFFSR_108 OR2X2_6/gnd DFFSR_92/S FILL
XDFFPOSX1_2 AOI21X1_1/A CLKBUF1_49/Y NOR2X1_59/Y DFFSR_1/gnd DFFSR_1/S DFFPOSX1
XFILL_4_DFFPOSX1_8 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_7_DFFPOSX1_22 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_34_DFFSR_212 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_5_AOI21X1_25 DFFSR_62/gnd DFFSR_208/S FILL
XAOI21X1_22 AOI21X1_22/A AOI21X1_22/B AOI21X1_22/C DFFSR_62/gnd OAI21X1_54/A DFFSR_62/S
+ AOI21X1
XFILL_10_DFFSR_111 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_4_AOI21X1_28 AND2X2_38/B DFFSR_23/S FILL
XFILL_24_DFFSR_215 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_52_4_1 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_50_DFFSR_50 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_39_DFFSR_90 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_3_AOI21X1_31 INVX1_39/gnd DFFSR_34/S FILL
XFILL_14_DFFSR_218 BUFX2_98/A DFFSR_32/S FILL
XFILL_2_AOI21X1_34 INVX1_39/gnd DFFSR_34/S FILL
XFILL_16_DFFPOSX1_41 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_50_6_2 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_6_DFFSR_47 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_5_NAND2X1_118 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_23_DFFSR_40 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_12_DFFSR_80 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_6_DFFSR_105 INVX1_1/gnd DFFSR_53/S FILL
XFILL_1_AOI21X1_37 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_0_NAND3X1_244 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_47_DFFSR_136 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_0_AOI21X1_40 INVX1_39/gnd DFFSR_54/S FILL
XFILL_37_DFFSR_139 DFFSR_34/gnd DFFSR_34/S FILL
XBUFX2_25 BUFX2_23/A BUFX2_8/gnd BUFX2_25/Y DFFSR_81/S BUFX2
XFILL_0_DFFSR_215 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_27_DFFSR_142 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_3_OAI21X1_100 INVX1_3/gnd DFFSR_79/S FILL
XFILL_26_DFFPOSX1_30 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_31_2 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_41_DFFSR_246 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_47_DFFSR_97 INVX1_1/gnd DFFSR_97/S FILL
XFILL_3_INVX1_189 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_17_DFFSR_145 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_8_OAI21X1_64 INVX1_1/gnd DFFSR_53/S FILL
XFILL_31_DFFSR_249 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_1_NAND3X1_178 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_8_AND2X2_6 BUFX2_99/A DFFSR_7/S FILL
XFILL_7_OAI21X1_67 INVX1_1/gnd DFFSR_97/S FILL
XFILL_6_NAND2X1_85 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_21_DFFSR_252 AND2X2_38/B DFFSR_23/S FILL
XFILL_3_INVX1_41 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_31_DFFSR_47 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_3_DFFSR_94 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_18_5_0 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_2_NOR2X1_24 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_20_DFFSR_87 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_5_NAND2X1_88 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_11_DFFSR_255 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_6_OAI21X1_70 INVX1_3/gnd DFFSR_23/S FILL
XNAND2X1_85 AND2X2_33/Y AND2X2_37/Y NOR3X1_6/gnd NAND2X1_85/Y DFFSR_91/S NAND2X1
XFILL_4_NAND2X1_91 INVX1_39/gnd DFFSR_54/S FILL
XFILL_5_OAI21X1_73 DFFSR_46/gnd DFFSR_54/S FILL
XOAI21X1_70 OR2X2_3/A OAI21X1_72/B AOI21X1_31/Y INVX1_3/gnd OAI21X1_70/Y DFFSR_23/S
+ OAI21X1
XFILL_2_NAND3X1_112 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_3_DFFSR_142 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_3_NAND2X1_94 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_4_OAI21X1_76 INVX1_1/gnd DFFSR_53/S FILL
XFILL_2_BUFX2_32 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_44_DFFSR_173 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_3_OAI21X1_79 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_2_NAND2X1_97 INVX1_1/gnd DFFSR_97/S FILL
XFILL_7_DFFSR_249 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_1_DFFSR_7 BUFX2_79/A DFFSR_7/S FILL
XFILL_4_NAND2X1_148 INVX1_67/gnd DFFSR_175/S FILL
XFILL_34_DFFSR_176 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_2_OAI21X1_82 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_48_DFFSR_280 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_24_DFFSR_179 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_50_DFFSR_14 INVX1_1/gnd DFFSR_53/S FILL
XFILL_1_OAI21X1_85 INVX1_39/gnd DFFSR_54/S FILL
XFILL_0_INVX1_88 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_28_DFFSR_94 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_39_DFFSR_54 INVX1_39/gnd DFFSR_54/S FILL
XFILL_14_DFFSR_182 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_0_OAI21X1_88 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_6_DFFSR_11 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_12_DFFSR_44 DFFSR_4/gnd DFFSR_98/S FILL
XBUFX2_3 BUFX2_3/A BUFX2_8/gnd BUFX2_3/Y DFFSR_81/S BUFX2
XFILL_1_OAI21X1_9 INVX1_67/gnd DFFSR_201/S FILL
XFILL_47_DFFSR_100 INVX1_1/gnd DFFSR_97/S FILL
XFILL_0_NAND3X1_208 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_37_DFFSR_103 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_0_DFFSR_179 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_27_DFFSR_106 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_41_DFFSR_210 BUFX2_98/A DFFSR_6/S FILL
XFILL_3_INVX1_153 INVX1_67/gnd DFFSR_175/S FILL
XFILL_47_DFFSR_61 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_6_AND2X2_20 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_17_DFFSR_109 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_8_OAI21X1_28 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_28_0_0 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_31_DFFSR_213 INVX1_3/gnd DFFSR_23/S FILL
XFILL_1_NAND3X1_142 INVX1_67/gnd DFFSR_175/S FILL
XFILL_6_NAND2X1_49 INVX1_3/gnd DFFSR_79/S FILL
XFILL_7_OAI21X1_31 AND2X2_38/B DFFSR_23/S FILL
XFILL_21_DFFSR_216 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_3_DFFSR_58 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_31_DFFSR_11 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_6_DFFPOSX1_16 INVX1_67/gnd DFFSR_175/S FILL
XFILL_20_DFFSR_51 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_6_OAI21X1_34 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_5_NAND2X1_52 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_11_DFFSR_219 INVX1_67/gnd DFFSR_175/S FILL
XFILL_3_NAND2X1_178 INVX1_1/gnd DFFSR_53/S FILL
XFILL_26_2_1 INVX1_3/gnd DFFSR_23/S FILL
XNAND2X1_49 DFFSR_239/Q NOR2X1_34/Y INVX1_3/gnd OAI21X1_15/C DFFSR_79/S NAND2X1
XFILL_5_OAI21X1_37 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_4_NAND2X1_55 INVX1_39/gnd DFFSR_34/S FILL
XFILL_8_1_0 XOR2X1_1/gnd DFFSR_151/S FILL
XOAI21X1_34 INVX1_147/A INVX1_149/Y INVX1_148/Y BUFX2_7/gnd AOI21X1_18/A DFFSR_151/S
+ OAI21X1
XFILL_3_DFFSR_106 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_3_NAND2X1_58 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_4_OAI21X1_40 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_24_4_2 AND2X2_38/B DFFSR_59/S FILL
XFILL_44_DFFSR_137 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_2_NAND2X1_61 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_3_OAI21X1_43 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_15_DFFPOSX1_35 INVX1_39/gnd DFFSR_54/S FILL
XFILL_46_DFFSR_7 BUFX2_79/A DFFSR_7/S FILL
XFILL_6_3_1 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_7_DFFSR_213 INVX1_3/gnd DFFSR_23/S FILL
XFILL_4_NAND2X1_112 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_34_DFFSR_140 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_1_NAND2X1_64 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_48_DFFSR_244 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_2_OAI21X1_46 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_11_AOI22X1_12 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_24_DFFSR_143 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_38_DFFSR_247 BUFX2_99/A DFFSR_7/S FILL
XFILL_0_NAND2X1_67 AND2X2_38/B DFFSR_59/S FILL
XFILL_1_OAI21X1_49 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_0_INVX1_190 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_28_DFFSR_58 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_0_INVX1_52 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_17_DFFSR_98 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_39_DFFSR_18 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_10_AOI22X1_15 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_4_5_2 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_14_DFFSR_146 BUFX2_79/A DFFSR_7/S FILL
XFILL_0_OAI21X1_52 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_28_DFFSR_250 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_53_2 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_25_DFFPOSX1_24 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_18_DFFSR_253 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_9_AOI22X1_18 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_1_INVX1_9 BUFX2_99/A DFFSR_7/S FILL
XFILL_8_AOI22X1_21 AND2X2_38/B DFFSR_59/S FILL
XFILL_0_NAND3X1_172 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_7_AOI22X1_24 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_5_DFFPOSX1_46 INVX1_39/gnd DFFSR_34/S FILL
XFILL_0_DFFSR_143 OR2X2_2/gnd DFFSR_216/S FILL
XDFFSR_253 BUFX2_94/A CLKBUF1_6/Y BUFX2_66/Y DFFSR_1/S INVX1_96/A DFFSR_34/gnd DFFSR_1/S
+ DFFSR
XFILL_6_AOI22X1_27 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_41_DFFSR_174 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_3_INVX1_117 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_47_DFFSR_25 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_36_DFFSR_65 BUFX2_79/A DFFSR_7/S FILL
XFILL_4_DFFSR_250 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_31_DFFSR_177 DFFSR_46/gnd DFFSR_54/S FILL
XAOI22X1_27 AOI22X1_28/A NAND2X1_98/Y AOI22X1_29/C INVX1_174/A OR2X2_6/gnd OAI21X1_69/B
+ DFFSR_92/S AOI22X1
XFILL_1_NAND3X1_106 INVX1_3/gnd DFFSR_23/S FILL
XFILL_6_NAND2X1_13 BUFX2_99/A DFFSR_92/S FILL
XFILL_21_DFFSR_180 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_3_DFFSR_22 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_20_DFFSR_15 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_5_NAND2X1_16 BUFX2_79/A DFFSR_7/S FILL
XFILL_11_DFFSR_183 INVX1_67/gnd DFFSR_175/S FILL
XFILL_3_NAND2X1_142 INVX1_67/gnd DFFSR_175/S FILL
XNAND2X1_13 DFFSR_114/D NOR2X1_5/Y BUFX2_99/A OAI21X1_2/C DFFSR_92/S NAND2X1
XFILL_4_NAND2X1_19 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_6_NOR2X1_59 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_8_OAI21X1_7 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_3_NAND2X1_22 BUFX2_99/A DFFSR_7/S FILL
XFILL_2_NOR2X1_3 XOR2X1_4/gnd DFFSR_91/S FILL
XDFFPOSX1_16 AOI21X1_7/C CLKBUF1_44/Y OAI21X1_28/Y INVX1_67/gnd DFFSR_175/S DFFPOSX1
XFILL_44_DFFSR_101 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_12_DFFSR_5 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_2_NAND2X1_25 BUFX2_99/A DFFSR_7/S FILL
XFILL_44_DFFSR_72 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_7_DFFSR_177 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_34_DFFSR_104 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_1_NAND2X1_28 AND2X2_38/B DFFSR_59/S FILL
XFILL_2_OAI21X1_10 BUFX2_79/A DFFSR_7/S FILL
XFILL_48_DFFSR_208 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_24_DFFSR_107 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_8_NAND3X1_84 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_38_DFFSR_211 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_0_NAND2X1_31 INVX1_3/gnd DFFSR_23/S FILL
XFILL_1_OAI21X1_13 INVX1_39/gnd DFFSR_54/S FILL
XFILL_28_DFFSR_22 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_0_DFFSR_69 BUFX2_98/A DFFSR_32/S FILL
XFILL_0_INVX1_16 BUFX2_99/A DFFSR_7/S FILL
XFILL_17_DFFSR_62 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_0_INVX1_154 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_3_AND2X2_21 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_14_DFFSR_110 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_7_NAND3X1_87 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_4_BUFX2_97 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_0_OAI21X1_16 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_28_DFFSR_214 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_6_NAND3X1_90 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_18_DFFSR_217 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_5_NAND3X1_93 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_0_NAND3X1_136 DFFSR_1/gnd DFFSR_81/S FILL
XNAND3X1_90 DFFSR_156/D AND2X2_18/B BUFX2_29/Y OR2X2_1/gnd AND2X2_22/B DFFSR_59/S
+ NAND3X1
XFILL_9_NAND3X1_191 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_4_NAND3X1_96 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_33_DFFSR_1 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_5_DFFPOSX1_10 INVX1_67/gnd DFFSR_201/S FILL
XFILL_3_NAND3X1_99 OR2X2_1/gnd DFFSR_51/S FILL
XDFFSR_217 DFFSR_217/Q CLKBUF1_34/Y BUFX2_62/Y DFFSR_201/S INVX1_64/A BUFX2_72/gnd
+ DFFSR_201/S DFFSR
XFILL_0_DFFSR_107 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_2_NAND2X1_172 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_41_DFFSR_138 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_36_DFFSR_29 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_8_DFFSR_76 BUFX2_79/A DFFSR_7/S FILL
XFILL_25_DFFSR_69 BUFX2_98/A DFFSR_32/S FILL
XFILL_4_DFFSR_214 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_31_DFFSR_141 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_45_DFFSR_245 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_7_CLKBUF1_9 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_21_DFFSR_144 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_14_DFFPOSX1_29 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_35_DFFSR_248 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_3_NAND2X1_106 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_11_DFFSR_147 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_25_DFFSR_251 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_6_NOR2X1_23 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_15_DFFSR_254 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_10_OAI22X1_27 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_44_DFFSR_36 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_33_DFFSR_76 BUFX2_79/A DFFSR_7/S FILL
XFILL_7_DFFSR_141 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_24_DFFPOSX1_18 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_48_DFFSR_172 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_8_NAND3X1_48 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_9_OAI22X1_30 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_38_DFFSR_175 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_0_DFFSR_33 BUFX2_98/A DFFSR_32/S FILL
XFILL_0_INVX1_118 BUFX2_98/A DFFSR_6/S FILL
XFILL_17_DFFSR_26 BUFX2_79/A DFFSR_6/S FILL
XFILL_8_NAND3X1_221 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_1_DFFSR_251 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_7_NAND3X1_51 BUFX2_99/A DFFSR_7/S FILL
XFILL_25_5_0 AND2X2_38/B DFFSR_23/S FILL
XFILL_4_BUFX2_61 AND2X2_38/B DFFSR_59/S FILL
XFILL_8_OAI22X1_33 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_28_DFFSR_178 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_4_DFFPOSX1_40 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_7_OAI22X1_36 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_6_NAND3X1_54 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_18_DFFSR_181 INVX1_3/gnd DFFSR_79/S FILL
XFILL_5_NAND3X1_57 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_6_OAI22X1_39 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_0_NAND3X1_100 AND2X2_38/B DFFSR_59/S FILL
XNAND3X1_54 DFFSR_79/D BUFX2_15/Y NOR2X1_2/Y OR2X2_3/gnd NAND3X1_55/B DFFSR_60/S NAND3X1
XFILL_4_NAND3X1_60 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_5_OAI22X1_42 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_41_DFFSR_83 INVX1_3/gnd DFFSR_79/S FILL
XFILL_5_6_0 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_3_NOR2X1_60 DFFSR_34/gnd DFFSR_34/S FILL
XOAI22X1_39 INVX1_94/Y OAI22X1_45/B INVX1_95/Y OAI22X1_45/D BUFX2_77/gnd NOR2X1_48/A
+ DFFSR_5/S OAI22X1
XFILL_4_OAI22X1_45 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_3_NAND3X1_63 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_5_OAI21X1_8 BUFX2_99/A DFFSR_7/S FILL
XFILL_2_NAND2X1_136 BUFX2_72/gnd DFFSR_276/S FILL
XDFFSR_181 INVX1_90/A CLKBUF1_12/Y BUFX2_70/Y DFFSR_79/S INVX1_91/A INVX1_3/gnd DFFSR_79/S
+ DFFSR
XFILL_2_NAND3X1_66 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_41_DFFSR_102 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_3_OAI22X1_48 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_8_DFFSR_40 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_25_DFFSR_33 BUFX2_98/A DFFSR_32/S FILL
XFILL_14_DFFSR_73 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_4_DFFSR_178 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_31_DFFSR_105 INVX1_1/gnd DFFSR_53/S FILL
XFILL_1_NAND3X1_69 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_2_OAI22X1_51 INVX1_39/gnd DFFSR_54/S FILL
XFILL_45_DFFSR_209 BUFX2_72/gnd DFFSR_276/S FILL
XNAND2X1_2 NOR2X1_1/Y BUFX2_11/Y BUFX2_99/A OAI22X1_7/B DFFSR_7/S NAND2X1
XFILL_21_DFFSR_108 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_0_NAND3X1_72 INVX1_39/gnd DFFSR_34/S FILL
XFILL_35_DFFSR_212 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_0_OAI21X1_118 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_23_DFFPOSX1_48 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_0_AND2X2_22 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_11_DFFSR_111 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_0_DFFSR_4 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_25_DFFSR_215 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_49_DFFSR_90 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_15_DFFSR_218 BUFX2_98/A DFFSR_32/S FILL
XOAI22X1_1 INVX1_1/Y OAI22X1_7/B INVX1_2/Y OAI22X1_7/D INVX1_1/gnd NOR2X1_3/B DFFSR_53/S
+ OAI22X1
XINVX1_74 INVX1_74/A BUFX2_99/A INVX1_74/Y DFFSR_92/S INVX1
XFILL_33_DFFSR_40 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_22_DFFSR_80 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_5_DFFSR_87 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_7_DFFSR_105 INVX1_1/gnd DFFSR_53/S FILL
XFILL_48_DFFSR_136 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_35_0_0 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_8_NAND3X1_12 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_38_DFFSR_139 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_8_NAND3X1_185 BUFX2_7/gnd DFFSR_216/S FILL
XINVX1_192 INVX1_192/A XOR2X1_1/gnd INVX1_192/Y DFFSR_151/S INVX1
XFILL_7_NAND3X1_15 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_4_BUFX2_25 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_1_DFFSR_215 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_18_4 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_28_DFFSR_142 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_33_2_1 INVX1_1/gnd DFFSR_53/S FILL
XFILL_1_NAND2X1_166 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_42_DFFSR_246 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_6_NAND3X1_18 BUFX2_79/A DFFSR_7/S FILL
XFILL_4_INVX1_189 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_18_DFFSR_145 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_32_DFFSR_249 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_24_DFFSR_8 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_5_NAND3X1_21 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_14_NOR3X1_4 NOR3X1_6/gnd DFFSR_91/S FILL
XNAND3X1_18 DFFSR_3/Q NOR2X1_4/Y BUFX2_16/Y BUFX2_79/A AND2X2_8/B DFFSR_7/S NAND3X1
XFILL_31_4_2 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_22_DFFSR_252 AND2X2_38/B DFFSR_23/S FILL
XFILL_4_NAND3X1_24 INVX1_1/gnd DFFSR_97/S FILL
XFILL_2_INVX1_81 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_30_DFFSR_87 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_41_DFFSR_47 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_3_NOR2X1_24 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_12_DFFSR_255 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_13_DFFPOSX1_23 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_3_NAND3X1_27 OR2X2_4/gnd DFFSR_3/S FILL
XDFFSR_145 INVX1_66/A CLKBUF1_25/Y BUFX2_67/Y DFFSR_201/S INVX1_67/A BUFX2_72/gnd
+ DFFSR_201/S DFFSR
XFILL_2_NAND2X1_100 INVX1_39/gnd DFFSR_54/S FILL
XFILL_3_OAI22X1_12 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_2_NAND3X1_30 BUFX2_79/A DFFSR_6/S FILL
XFILL_14_DFFSR_37 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_4_DFFSR_142 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_1_BUFX2_72 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_2_OAI22X1_15 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_1_NAND3X1_33 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_45_DFFSR_173 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_8_DFFSR_249 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_1_OAI22X1_18 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_0_NAND3X1_36 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_35_DFFSR_176 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_49_DFFSR_280 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_23_DFFPOSX1_12 AND2X2_38/B DFFSR_23/S FILL
XFILL_0_OAI22X1_21 BUFX2_98/A DFFSR_32/S FILL
XFILL_45_DFFSR_4 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_25_DFFSR_179 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_38_DFFSR_94 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_49_DFFSR_54 INVX1_39/gnd DFFSR_54/S FILL
XFILL_7_NAND3X1_215 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_15_DFFSR_182 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_3_DFFPOSX1_34 OR2X2_2/gnd DFFSR_216/S FILL
XDFFSR_91 DFFSR_91/Q DFFSR_83/CLK DFFSR_73/R DFFSR_91/S DFFSR_83/Q XOR2X1_4/gnd DFFSR_91/S
+ DFFSR
XINVX1_38 DFFSR_54/Q AND2X2_38/B INVX1_38/Y DFFSR_23/S INVX1
XFILL_22_DFFSR_44 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_5_DFFSR_51 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_11_DFFSR_84 BUFX2_99/A DFFSR_7/S FILL
XFILL_0_NOR2X1_61 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_2_OAI21X1_9 INVX1_67/gnd DFFSR_201/S FILL
XFILL_48_DFFSR_100 INVX1_1/gnd DFFSR_97/S FILL
XFILL_38_DFFSR_103 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_8_NAND3X1_149 DFFSR_1/gnd DFFSR_1/S FILL
XINVX1_156 INVX1_156/A DFFSR_62/gnd INVX1_156/Y DFFSR_62/S INVX1
XFILL_1_DFFSR_179 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_0_INVX1_6 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_28_DFFSR_106 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_42_DFFSR_210 BUFX2_98/A DFFSR_6/S FILL
XFILL_1_NAND2X1_130 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_4_INVX1_153 INVX1_67/gnd DFFSR_175/S FILL
XFILL_7_AND2X2_20 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_18_DFFSR_109 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_32_DFFSR_213 INVX1_3/gnd DFFSR_23/S FILL
XFILL_22_DFFSR_216 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_2_INVX1_45 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_41_DFFSR_11 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_2_DFFSR_98 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_19_DFFSR_91 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_30_DFFSR_51 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_12_DFFSR_219 INVX1_67/gnd DFFSR_175/S FILL
XDFFSR_109 DFFSR_109/Q DFFSR_93/CLK DFFSR_5/R DFFSR_4/S AOI22X1_5/B DFFSR_4/gnd DFFSR_4/S
+ DFFSR
XFILL_22_DFFPOSX1_42 INVX1_39/gnd DFFSR_34/S FILL
XFILL_4_DFFSR_106 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_1_BUFX2_36 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_6_NAND3X1_245 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_45_DFFSR_137 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_8_DFFSR_213 INVX1_3/gnd DFFSR_23/S FILL
XFILL_35_DFFSR_140 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_49_DFFSR_244 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_11_DFFSR_2 BUFX2_79/A DFFSR_7/S FILL
XFILL_25_DFFSR_143 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_1_INVX1_190 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_38_DFFSR_58 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_39_DFFSR_247 BUFX2_99/A DFFSR_7/S FILL
XFILL_49_DFFSR_18 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_27_DFFSR_98 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_15_DFFSR_146 BUFX2_79/A DFFSR_7/S FILL
XFILL_7_NAND3X1_179 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_29_DFFSR_250 DFFSR_8/gnd DFFSR_8/S FILL
XDFFSR_55 DFFSR_15/D CLKBUF1_37/Y DFFSR_15/R DFFSR_4/S DFFSR_55/D DFFSR_4/gnd DFFSR_4/S
+ DFFSR
XFILL_0_NAND2X1_160 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_19_DFFSR_253 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_5_DFFSR_15 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_11_DFFSR_48 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_0_NOR2X1_25 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_8_NAND3X1_113 DFFSR_62/gnd DFFSR_208/S FILL
XINVX1_120 INVX1_120/A DFFSR_62/gnd INVX1_120/Y DFFSR_208/S INVX1
XFILL_1_DFFSR_143 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_12_DFFPOSX1_17 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_42_DFFSR_174 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_4_INVX1_117 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_46_DFFSR_65 BUFX2_79/A DFFSR_7/S FILL
XFILL_5_DFFSR_250 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_32_DFFSR_177 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_22_DFFSR_180 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_30_DFFSR_15 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_19_DFFSR_55 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_2_DFFSR_62 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_12_DFFSR_183 INVX1_67/gnd DFFSR_175/S FILL
XFILL_6_BUFX2_90 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_9_OAI21X1_7 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_20_CLKBUF1_45 BUFX2_79/A DFFSR_7/S FILL
XFILL_6_NAND3X1_209 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_45_DFFSR_101 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_32_5_0 INVX1_1/gnd DFFSR_97/S FILL
XFILL_2_DFFPOSX1_28 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_19_CLKBUF1_48 INVX1_3/gnd DFFSR_79/S FILL
XFILL_8_DFFSR_177 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_35_DFFSR_104 DFFSR_28/gnd DFFSR_8/S FILL
XAND2X2_24 AND2X2_24/A AND2X2_24/B BUFX2_8/gnd AND2X2_24/Y DFFSR_51/S AND2X2
XFILL_49_DFFSR_208 DFFSR_62/gnd DFFSR_208/S FILL
XNAND3X1_245 INVX1_170/A AOI21X1_44/B OR2X2_4/Y OR2X2_4/gnd NAND3X1_245/Y DFFSR_3/S
+ NAND3X1
XFILL_25_DFFSR_107 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_39_DFFSR_211 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_38_DFFSR_22 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_1_INVX1_154 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_4_AND2X2_21 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_27_DFFSR_62 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_15_DFFSR_110 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_7_NAND3X1_143 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_29_DFFSR_214 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_11_DFFPOSX1_47 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_19_DFFSR_217 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_0_NAND2X1_124 OR2X2_2/gnd DFFSR_216/S FILL
XDFFSR_19 INVX1_21/A CLKBUF1_7/Y DFFSR_3/R DFFSR_8/S INVX1_22/A DFFSR_28/gnd DFFSR_8/S
+ DFFSR
XFILL_11_DFFSR_12 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_1_DFFSR_107 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_21_DFFPOSX1_36 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_42_DFFSR_138 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_46_DFFSR_29 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_35_DFFSR_69 BUFX2_98/A DFFSR_32/S FILL
XFILL_5_DFFSR_214 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_32_DFFSR_141 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_46_DFFSR_245 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_5_NAND3X1_239 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_8_CLKBUF1_9 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_22_DFFSR_144 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_2_DFFSR_26 BUFX2_79/A DFFSR_6/S FILL
XFILL_36_DFFSR_248 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_19_DFFSR_19 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_6_BUFX2_54 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_12_DFFSR_147 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_26_DFFSR_251 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_42_0_0 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_16_DFFSR_254 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_1_NOR2X1_7 BUFX2_98/A DFFSR_32/S FILL
XFILL_6_NAND3X1_173 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_43_DFFSR_76 BUFX2_79/A DFFSR_7/S FILL
XFILL_19_CLKBUF1_12 AND2X2_38/B DFFSR_23/S FILL
XFILL_40_2_1 BUFX2_98/A DFFSR_6/S FILL
XFILL_8_DFFSR_141 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_18_CLKBUF1_15 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_49_DFFSR_172 DFFSR_46/gnd DFFSR_62/S FILL
XNAND3X1_209 AOI21X1_22/A OAI21X1_58/C AOI21X1_22/B DFFSR_46/gnd AOI21X1_32/B DFFSR_62/S
+ NAND3X1
XFILL_39_DFFSR_175 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_17_CLKBUF1_18 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_1_INVX1_118 BUFX2_98/A DFFSR_6/S FILL
XFILL_27_DFFSR_26 BUFX2_79/A DFFSR_6/S FILL
XFILL_16_DFFSR_66 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_0_BUFX2_100 BUFX2_79/A DFFSR_6/S FILL
XFILL_38_4_2 BUFX2_79/A DFFSR_7/S FILL
XFILL_2_DFFSR_251 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_7_NAND3X1_107 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_16_CLKBUF1_21 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_29_DFFSR_178 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_11_DFFPOSX1_11 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_15_CLKBUF1_24 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_19_DFFSR_181 INVX1_3/gnd DFFSR_79/S FILL
XNOR2X1_63 AND2X2_28/Y NOR2X1_63/B INVX1_3/gnd NOR2X1_63/Y DFFSR_23/S NOR2X1
XFILL_14_CLKBUF1_27 INVX1_1/gnd DFFSR_97/S FILL
XFILL_3_XOR2X1_3 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_51_DFFSR_83 INVX1_3/gnd DFFSR_79/S FILL
XFILL_23_DFFSR_5 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_13_CLKBUF1_30 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_4_NOR2X1_60 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_6_OAI21X1_8 BUFX2_99/A DFFSR_7/S FILL
XFILL_12_CLKBUF1_33 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_42_DFFSR_102 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_7_DFFSR_80 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_35_DFFSR_33 BUFX2_98/A DFFSR_32/S FILL
XFILL_11_CLKBUF1_36 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_24_DFFSR_73 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_5_DFFSR_178 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_32_DFFSR_105 INVX1_1/gnd DFFSR_53/S FILL
XFILL_46_DFFSR_209 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_10_CLKBUF1_39 INVX1_1/gnd DFFSR_53/S FILL
XFILL_5_NAND3X1_203 INVX1_1/gnd DFFSR_97/S FILL
XFILL_22_DFFSR_108 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_36_DFFSR_212 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_1_DFFPOSX1_22 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_1_AND2X2_22 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_12_DFFSR_111 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_6_BUFX2_18 BUFX2_98/A DFFSR_32/S FILL
XFILL_9_CLKBUF1_42 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_26_DFFSR_215 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_16_DFFSR_218 BUFX2_98/A DFFSR_32/S FILL
XFILL_8_CLKBUF1_45 BUFX2_79/A DFFSR_7/S FILL
XFILL_44_DFFSR_1 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_6_NAND3X1_137 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_7_CLKBUF1_48 INVX1_3/gnd DFFSR_79/S FILL
XFILL_10_DFFPOSX1_41 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_43_DFFSR_40 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_4_INVX1_74 BUFX2_99/A DFFSR_92/S FILL
XFILL_32_DFFSR_80 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_8_DFFSR_105 INVX1_1/gnd DFFSR_53/S FILL
XFILL_49_DFFSR_136 NOR3X1_6/gnd DFFSR_79/S FILL
XNAND3X1_173 INVX1_160/Y AOI21X1_30/B NAND2X1_85/Y XOR2X1_4/gnd AOI21X1_28/A DFFSR_91/S
+ NAND3X1
XFILL_39_DFFSR_139 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_16_DFFSR_30 BUFX2_98/A DFFSR_32/S FILL
XFILL_22_1 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_2_DFFSR_215 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_3_BUFX2_65 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_29_DFFSR_142 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_43_DFFSR_246 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_20_DFFPOSX1_30 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_19_DFFSR_145 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_33_DFFSR_249 BUFX2_72/gnd DFFSR_276/S FILL
XNOR2X1_27 NOR2X1_27/A NOR2X1_27/B DFFSR_8/gnd NOR2X1_27/Y DFFSR_60/S NOR2X1
XFILL_4_NAND3X1_233 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_23_DFFSR_252 AND2X2_38/B DFFSR_23/S FILL
XFILL_40_DFFSR_87 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_4_NOR2X1_24 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_13_DFFSR_255 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_24_DFFSR_37 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_7_DFFSR_44 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_13_DFFSR_77 BUFX2_98/A DFFSR_32/S FILL
XFILL_5_DFFSR_142 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_14_0_1 INVX1_39/gnd DFFSR_54/S FILL
XFILL_46_DFFSR_173 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_5_NAND3X1_167 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_9_DFFSR_249 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_36_DFFSR_176 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_50_DFFSR_280 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_26_DFFSR_179 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_12_2_2 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_48_DFFSR_94 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_16_DFFSR_182 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_6_NAND3X1_101 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_7_CLKBUF1_12 AND2X2_38/B DFFSR_23/S FILL
XFILL_4_DFFSR_91 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_4_INVX1_38 AND2X2_38/B DFFSR_23/S FILL
XFILL_32_DFFSR_44 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_21_DFFSR_84 BUFX2_99/A DFFSR_7/S FILL
XFILL_1_NOR2X1_61 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_6_CLKBUF1_15 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_3_OAI21X1_9 INVX1_67/gnd DFFSR_201/S FILL
XFILL_49_DFFSR_100 INVX1_1/gnd DFFSR_97/S FILL
XFILL_5_CLKBUF1_18 OR2X2_1/gnd DFFSR_51/S FILL
XNAND3X1_137 BUFX2_58/Y INVX1_133/A NAND2X1_59/A BUFX2_7/gnd INVX1_136/A DFFSR_216/S
+ NAND3X1
XFILL_39_DFFSR_103 DFFSR_8/gnd DFFSR_60/S FILL
XCLKBUF1_15 BUFX2_3/Y DFFSR_46/gnd CLKBUF1_15/Y DFFSR_62/S CLKBUF1
XFILL_5_5 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_4_CLKBUF1_21 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_2_DFFSR_179 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_3_BUFX2_29 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_29_DFFSR_106 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_43_DFFSR_210 BUFX2_98/A DFFSR_6/S FILL
XFILL_3_CLKBUF1_24 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_8_AND2X2_20 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_19_DFFSR_109 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_6_OAI21X1_119 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_2_CLKBUF1_27 INVX1_1/gnd DFFSR_97/S FILL
XFILL_33_DFFSR_213 INVX1_3/gnd DFFSR_23/S FILL
XFILL_23_DFFSR_216 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_1_CLKBUF1_30 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_4_NAND3X1_197 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_39_5_0 BUFX2_79/A DFFSR_6/S FILL
XFILL_29_DFFSR_91 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_40_DFFSR_51 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_51_DFFSR_11 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_1_INVX1_85 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_13_DFFSR_219 INVX1_67/gnd DFFSR_175/S FILL
XFILL_0_DFFPOSX1_16 INVX1_67/gnd DFFSR_175/S FILL
XFILL_0_CLKBUF1_33 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_13_DFFSR_41 BUFX2_98/A DFFSR_6/S FILL
XFILL_5_DFFSR_106 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_0_BUFX2_76 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_46_DFFSR_137 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_5_NAND3X1_131 AND2X2_38/B DFFSR_59/S FILL
XFILL_9_DFFSR_213 INVX1_3/gnd DFFSR_23/S FILL
XFILL_36_DFFSR_140 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_50_DFFSR_244 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_26_DFFSR_143 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_35_DFFSR_8 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_2_INVX1_190 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_48_DFFSR_58 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_40_DFFSR_247 BUFX2_99/A DFFSR_7/S FILL
XFILL_37_DFFSR_98 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_16_DFFSR_146 BUFX2_79/A DFFSR_7/S FILL
XFILL_44_1 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_30_DFFSR_250 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_20_DFFSR_253 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_4_DFFSR_55 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_21_DFFSR_48 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_10_DFFSR_88 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_19_DFFPOSX1_24 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_1_NOR2X1_25 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_10_DFFSR_256 DFFSR_8/gnd DFFSR_60/S FILL
XNAND3X1_101 DFFSR_141/Q BUFX2_33/Y BUFX2_26/Y XOR2X1_4/gnd NAND3X1_103/A DFFSR_91/S
+ NAND3X1
XFILL_3_NAND3X1_227 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_2_DFFSR_143 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_43_DFFSR_174 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_6_DFFSR_250 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_49_0_0 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_33_DFFSR_177 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_4_NAND3X1_161 AND2X2_38/B DFFSR_23/S FILL
XFILL_23_DFFSR_180 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_40_DFFSR_15 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_29_DFFSR_55 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_1_INVX1_49 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_18_DFFSR_95 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_13_DFFSR_183 INVX1_67/gnd DFFSR_175/S FILL
XFILL_47_2_1 DFFSR_8/gnd DFFSR_60/S FILL
XOAI21X1_119 OR2X2_6/B OR2X2_6/A XOR2X1_15/Y OR2X2_6/gnd AOI21X1_71/A DFFSR_53/S OAI21X1
XFILL_9_DFFPOSX1_35 INVX1_39/gnd DFFSR_54/S FILL
XFILL_45_4_2 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_0_BUFX2_40 INVX1_1/gnd DFFSR_97/S FILL
XFILL_46_DFFSR_101 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_9_DFFSR_177 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_36_DFFSR_104 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_50_DFFSR_208 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_26_DFFSR_107 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_40_DFFSR_211 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_48_DFFSR_22 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_2_INVX1_154 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_5_AND2X2_21 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_37_DFFSR_62 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_16_DFFSR_110 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_30_DFFSR_214 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_20_DFFSR_217 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_4_DFFSR_19 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_21_DFFSR_12 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_10_DFFSR_52 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_5_OAI21X1_113 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_10_DFFSR_220 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_13_3_0 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_3_NAND3X1_191 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_2_DFFSR_107 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_22_DFFSR_2 BUFX2_79/A DFFSR_7/S FILL
XFILL_43_DFFSR_138 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_11_5_1 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_45_DFFSR_69 BUFX2_98/A DFFSR_32/S FILL
XFILL_6_DFFSR_214 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_33_DFFSR_141 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_47_DFFSR_245 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_9_CLKBUF1_9 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_4_NAND3X1_125 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_23_DFFSR_144 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_37_DFFSR_248 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_29_DFFSR_19 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_1_INVX1_13 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_1_DFFSR_66 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_18_DFFSR_59 AND2X2_38/B DFFSR_59/S FILL
XFILL_13_DFFSR_147 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_5_BUFX2_94 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_6_BUFX2_3 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_27_DFFSR_251 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_6_NAND2X1_161 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_49_6 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_17_DFFSR_254 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_9_DFFSR_141 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_18_DFFPOSX1_18 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_50_DFFSR_172 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_40_DFFSR_175 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_2_INVX1_118 BUFX2_98/A DFFSR_6/S FILL
XFILL_9_DFFSR_73 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_26_DFFSR_66 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_1_BUFX2_100 BUFX2_79/A DFFSR_6/S FILL
XFILL_37_DFFSR_26 BUFX2_79/A DFFSR_6/S FILL
XFILL_3_DFFSR_251 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_18_DFFPOSX1_3 INVX1_39/gnd DFFSR_34/S FILL
XFILL_2_NAND3X1_221 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_30_DFFSR_178 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_17_DFFPOSX1_6 AND2X2_38/B DFFSR_23/S FILL
XFILL_20_DFFSR_181 INVX1_3/gnd DFFSR_79/S FILL
XFILL_10_DFFSR_16 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_16_DFFPOSX1_9 INVX1_67/gnd DFFSR_201/S FILL
XFILL_10_DFFSR_184 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_21_0_1 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_3_NAND3X1_155 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_5_NOR2X1_60 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_7_OAI21X1_8 BUFX2_99/A DFFSR_7/S FILL
XFILL_8_DFFPOSX1_29 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_43_DFFSR_102 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_45_DFFSR_33 BUFX2_98/A DFFSR_32/S FILL
XFILL_34_DFFSR_73 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_6_DFFSR_178 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_19_2_2 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_33_DFFSR_105 INVX1_1/gnd DFFSR_53/S FILL
XFILL_47_DFFSR_209 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_1_1_1 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_23_DFFSR_108 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_37_DFFSR_212 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_1_DFFSR_30 BUFX2_98/A DFFSR_32/S FILL
XFILL_18_DFFSR_23 AND2X2_38/B DFFSR_23/S FILL
XFILL_2_AND2X2_22 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_13_DFFSR_111 DFFSR_8/gnd DFFSR_8/S FILL
XBUFX2_98 BUFX2_98/A BUFX2_79/A BUFX2_98/Y DFFSR_7/S BUFX2
XFILL_17_DFFPOSX1_48 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_5_BUFX2_58 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_10_OAI22X1_4 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_27_DFFSR_215 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_6_NAND2X1_125 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_17_DFFSR_218 BUFX2_98/A DFFSR_32/S FILL
XFILL_9_NOR3X1_4 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_9_AOI21X1_50 INVX1_67/gnd DFFSR_175/S FILL
XFILL_42_DFFSR_80 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_9_DFFSR_105 INVX1_1/gnd DFFSR_53/S FILL
XNAND2X1_161 DFFSR_201/S DFFPOSX1_29/Q BUFX2_72/gnd AOI21X1_56/B DFFSR_201/S NAND2X1
XFILL_50_DFFSR_136 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_8_AOI21X1_53 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_4_OAI21X1_107 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_27_DFFPOSX1_37 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_9_DFFSR_37 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_40_DFFSR_139 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_15_DFFSR_70 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_26_DFFSR_30 BUFX2_98/A DFFSR_32/S FILL
XFILL_7_AOI21X1_56 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_2_NAND3X1_185 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_3_DFFSR_215 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_30_DFFSR_142 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_46_5_0 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_6_AOI21X1_59 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_44_DFFSR_246 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_20_DFFSR_145 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_5_AOI21X1_62 INVX1_3/gnd DFFSR_23/S FILL
XFILL_34_DFFSR_249 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_10_DFFSR_148 INVX1_67/gnd DFFSR_175/S FILL
XAOI21X1_59 AOI21X1_59/A AOI21X1_59/B BUFX2_35/Y OR2X2_1/gnd AOI21X1_59/Y DFFSR_51/S
+ AOI21X1
XFILL_2_XOR2X1_7 BUFX2_98/A DFFSR_6/S FILL
XFILL_4_AOI21X1_65 INVX1_3/gnd DFFSR_23/S FILL
XFILL_24_DFFSR_252 AND2X2_38/B DFFSR_23/S FILL
XFILL_50_DFFSR_87 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_5_NOR2X1_24 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_13_DFFSR_9 BUFX2_79/A DFFSR_6/S FILL
XFILL_3_NAND3X1_119 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_3_AOI21X1_68 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_14_DFFSR_255 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_2_AOI21X1_71 BUFX2_99/A DFFSR_92/S FILL
XFILL_34_DFFSR_37 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_5_NAND2X1_155 BUFX2_79/A DFFSR_7/S FILL
XFILL_6_DFFSR_84 BUFX2_99/A DFFSR_7/S FILL
XFILL_6_DFFSR_142 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_23_DFFSR_77 BUFX2_98/A DFFSR_32/S FILL
XFILL_47_DFFSR_173 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_37_DFFSR_176 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_8_OR2X2_1 OR2X2_1/gnd DFFSR_59/S FILL
XBUFX2_62 BUFX2_60/A DFFSR_46/gnd BUFX2_62/Y DFFSR_62/S BUFX2
XFILL_5_BUFX2_22 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_17_DFFPOSX1_12 AND2X2_38/B DFFSR_23/S FILL
XFILL_0_DFFSR_252 AND2X2_38/B DFFSR_23/S FILL
XFILL_27_DFFSR_179 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_9_OAI21X1_98 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_17_DFFSR_182 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_34_DFFSR_5 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_15_NOR3X1_1 INVX1_3/gnd DFFSR_79/S FILL
XFILL_1_NAND3X1_215 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_42_DFFSR_44 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_31_DFFSR_84 BUFX2_99/A DFFSR_7/S FILL
XFILL_3_INVX1_78 DFFSR_46/gnd DFFSR_62/S FILL
XNAND2X1_125 BUFX2_54/Y INVX1_137/A OR2X2_2/gnd OAI21X1_94/C DFFSR_175/S NAND2X1
XFILL_2_NOR2X1_61 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_50_DFFSR_100 INVX1_1/gnd DFFSR_97/S FILL
XFILL_4_OAI21X1_9 INVX1_67/gnd DFFSR_201/S FILL
XFILL_8_AOI21X1_17 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_40_DFFSR_103 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_6_DFFPOSX1_3 INVX1_39/gnd DFFSR_34/S FILL
XFILL_9_2 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_7_AOI21X1_20 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_15_DFFSR_34 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_3_DFFSR_179 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_2_NAND3X1_149 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_2_BUFX2_69 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_30_DFFSR_106 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_5_DFFPOSX1_6 AND2X2_38/B DFFSR_23/S FILL
XFILL_6_AOI21X1_23 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_54_2_1 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_44_DFFSR_210 BUFX2_98/A DFFSR_6/S FILL
XFILL_9_AND2X2_20 OR2X2_6/gnd DFFSR_53/S FILL
XDFFPOSX1_3 AOI21X1_1/B CLKBUF1_49/Y AOI21X1_1/Y INVX1_39/gnd DFFSR_34/S DFFPOSX1
XFILL_20_DFFSR_109 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_7_DFFPOSX1_23 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_4_DFFPOSX1_9 INVX1_67/gnd DFFSR_201/S FILL
XFILL_5_AOI21X1_26 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_34_DFFSR_213 INVX1_3/gnd DFFSR_23/S FILL
XFILL_10_DFFSR_112 OR2X2_4/gnd DFFSR_32/S FILL
XAOI21X1_23 OAI21X1_43/Y NAND2X1_80/Y INVX1_156/Y DFFSR_62/gnd AOI21X1_23/Y DFFSR_62/S
+ AOI21X1
XFILL_4_AOI21X1_29 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_24_DFFSR_216 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_52_4_2 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_39_DFFSR_91 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_50_DFFSR_51 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_14_DFFSR_219 INVX1_67/gnd DFFSR_175/S FILL
XFILL_3_AOI21X1_32 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_16_DFFPOSX1_42 INVX1_39/gnd DFFSR_34/S FILL
XFILL_2_AOI21X1_35 INVX1_39/gnd DFFSR_54/S FILL
XFILL_6_DFFSR_48 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_5_NAND2X1_119 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_1_AOI21X1_38 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_23_DFFSR_41 BUFX2_98/A DFFSR_6/S FILL
XFILL_6_DFFSR_106 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_12_DFFSR_81 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_47_DFFSR_137 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_0_NAND3X1_245 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_0_AOI21X1_41 INVX1_39/gnd DFFSR_34/S FILL
XFILL_37_DFFSR_140 DFFSR_62/gnd DFFSR_208/S FILL
XBUFX2_26 BUFX2_23/A BUFX2_8/gnd BUFX2_26/Y DFFSR_51/S BUFX2
XFILL_0_DFFSR_216 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_27_DFFSR_143 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_3_OAI21X1_101 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_3_INVX1_190 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_41_DFFSR_247 BUFX2_99/A DFFSR_7/S FILL
XFILL_26_DFFPOSX1_31 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_31_3 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_47_DFFSR_98 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_20_3_0 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_17_DFFSR_146 BUFX2_79/A DFFSR_7/S FILL
XFILL_31_DFFSR_250 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_8_OAI21X1_65 INVX1_1/gnd DFFSR_53/S FILL
XFILL_1_NAND3X1_179 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_8_AND2X2_7 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_7_OAI21X1_68 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_6_NAND2X1_86 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_21_DFFSR_253 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_31_DFFSR_48 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_20_DFFSR_88 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_3_DFFSR_95 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_3_INVX1_42 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_18_5_1 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_2_NOR2X1_25 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_6_OAI21X1_71 INVX1_3/gnd DFFSR_79/S FILL
XFILL_5_NAND2X1_89 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_11_DFFSR_256 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_0_4_0 BUFX2_72/gnd DFFSR_276/S FILL
XNAND2X1_86 INVX1_135/A AND2X2_33/B NOR3X1_6/gnd NOR2X1_70/A DFFSR_91/S NAND2X1
XFILL_4_NAND2X1_92 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_5_OAI21X1_74 DFFSR_46/gnd DFFSR_62/S FILL
XOAI21X1_71 OAI21X1_69/A OAI21X1_69/B AOI21X1_31/Y INVX1_3/gnd OAI21X1_71/Y DFFSR_79/S
+ OAI21X1
XFILL_3_DFFSR_143 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_2_NAND3X1_113 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_4_OAI21X1_77 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_3_NAND2X1_95 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_2_BUFX2_33 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_44_DFFSR_174 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_3_OAI21X1_80 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_2_NAND2X1_98 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_7_DFFSR_250 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_1_DFFSR_8 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_4_NAND2X1_149 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_34_DFFSR_177 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_2_OAI21X1_83 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_24_DFFSR_180 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_50_DFFSR_15 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_39_DFFSR_55 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_1_OAI21X1_86 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_0_INVX1_89 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_28_DFFSR_95 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_14_DFFSR_183 INVX1_67/gnd DFFSR_175/S FILL
XFILL_0_OAI21X1_89 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_6_DFFSR_12 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_12_DFFSR_45 DFFSR_8/gnd DFFSR_60/S FILL
XBUFX2_4 BUFX2_3/A OR2X2_6/gnd BUFX2_4/Y DFFSR_92/S BUFX2
XFILL_47_DFFSR_101 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_0_NAND3X1_209 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_37_DFFSR_104 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_0_DFFSR_180 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_51_DFFSR_208 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_27_DFFSR_107 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_9_OAI21X1_26 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_41_DFFSR_211 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_3_INVX1_154 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_6_AND2X2_21 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_47_DFFSR_62 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_17_DFFSR_110 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_31_DFFSR_214 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_8_OAI21X1_29 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_28_0_1 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_1_NAND3X1_143 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_0_NAND2X1_1 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_21_DFFSR_217 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_7_OAI21X1_32 AND2X2_38/B DFFSR_59/S FILL
XFILL_6_NAND2X1_50 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_31_DFFSR_12 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_20_DFFSR_52 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_3_DFFSR_59 AND2X2_38/B DFFSR_59/S FILL
XFILL_6_DFFPOSX1_17 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_6_OAI21X1_35 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_3_NAND2X1_179 INVX1_1/gnd DFFSR_97/S FILL
XFILL_5_NAND2X1_53 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_11_DFFSR_220 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_26_2_2 INVX1_3/gnd DFFSR_23/S FILL
XNAND2X1_50 DFFSR_175/D AND2X2_18/Y DFFSR_62/gnd NAND2X1_50/Y DFFSR_62/S NAND2X1
XFILL_4_NAND2X1_56 AND2X2_38/B DFFSR_59/S FILL
XFILL_5_OAI21X1_38 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_8_1_1 XOR2X1_1/gnd DFFSR_151/S FILL
XOAI21X1_35 BUFX2_53/Y XOR2X1_3/Y OAI21X1_35/C BUFX2_7/gnd OAI21X1_35/Y DFFSR_216/S
+ OAI21X1
XFILL_3_DFFSR_107 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_4_OAI21X1_41 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_3_NAND2X1_59 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_44_DFFSR_138 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_15_DFFPOSX1_36 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_46_DFFSR_8 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_2_NAND2X1_62 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_3_OAI21X1_44 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_7_DFFSR_214 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_6_3_2 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_4_NAND2X1_113 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_34_DFFSR_141 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_2_OAI21X1_47 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_1_NAND2X1_65 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_48_DFFSR_245 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_24_DFFSR_144 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_1_OAI21X1_50 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_0_NAND2X1_68 AND2X2_38/B DFFSR_23/S FILL
XFILL_0_INVX1_191 INVX1_67/gnd DFFSR_175/S FILL
XFILL_38_DFFSR_248 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_39_DFFSR_19 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_0_INVX1_53 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_10_AOI22X1_16 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_17_DFFSR_99 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_28_DFFSR_59 AND2X2_38/B DFFSR_59/S FILL
XFILL_14_DFFSR_147 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_28_DFFSR_251 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_0_OAI21X1_53 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_53_3 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_25_DFFPOSX1_25 BUFX2_79/A DFFSR_6/S FILL
XFILL_9_AOI22X1_19 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_18_DFFSR_254 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_0_NAND3X1_173 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_8_AOI22X1_22 INVX1_3/gnd DFFSR_79/S FILL
XFILL_53_5_0 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_7_AOI22X1_25 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_5_DFFPOSX1_47 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_0_DFFSR_144 DFFSR_46/gnd DFFSR_62/S FILL
XDFFSR_254 BUFX2_95/A CLKBUF1_17/Y BUFX2_69/Y DFFSR_1/S DFFSR_246/Q DFFSR_34/gnd DFFSR_1/S
+ DFFSR
XFILL_6_AOI22X1_28 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_41_DFFSR_175 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_3_INVX1_118 BUFX2_98/A DFFSR_6/S FILL
XFILL_36_DFFSR_66 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_2_BUFX2_100 BUFX2_79/A DFFSR_6/S FILL
XFILL_47_DFFSR_26 BUFX2_79/A DFFSR_6/S FILL
XFILL_4_DFFSR_251 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_31_DFFSR_178 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_1_NAND3X1_107 BUFX2_8/gnd DFFSR_81/S FILL
XAOI22X1_28 AOI22X1_28/A NAND2X1_98/Y AOI22X1_26/C AOI22X1_26/D OR2X2_6/gnd OR2X2_3/A
+ DFFSR_53/S AOI22X1
XFILL_6_NAND2X1_14 BUFX2_98/A DFFSR_32/S FILL
XFILL_21_DFFSR_181 INVX1_3/gnd DFFSR_79/S FILL
XFILL_20_DFFSR_16 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_3_DFFSR_23 AND2X2_38/B DFFSR_23/S FILL
XFILL_3_NAND2X1_143 INVX1_67/gnd DFFSR_201/S FILL
XFILL_5_NAND2X1_17 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_11_DFFSR_184 OR2X2_1/gnd DFFSR_51/S FILL
XNAND2X1_14 DFFSR_34/Q AND2X2_5/Y BUFX2_98/A NAND2X1_14/Y DFFSR_32/S NAND2X1
XFILL_4_NAND2X1_20 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_6_NOR2X1_60 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_3_NAND2X1_23 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_8_OAI21X1_8 BUFX2_99/A DFFSR_7/S FILL
XFILL_2_NOR2X1_4 INVX1_1/gnd DFFSR_53/S FILL
XDFFPOSX1_17 INVX1_148/A CLKBUF1_48/Y OAI21X1_35/Y BUFX2_8/gnd DFFSR_51/S DFFPOSX1
XFILL_44_DFFSR_102 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_12_DFFSR_6 BUFX2_79/A DFFSR_6/S FILL
XFILL_2_NAND2X1_26 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_7_DFFSR_178 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_44_DFFSR_73 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_34_DFFSR_105 INVX1_1/gnd DFFSR_53/S FILL
XFILL_9_NAND3X1_82 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_1_NAND2X1_29 INVX1_3/gnd DFFSR_23/S FILL
XFILL_2_OAI21X1_11 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_48_DFFSR_209 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_24_DFFSR_108 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_8_NAND3X1_85 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_0_NAND2X1_32 INVX1_3/gnd DFFSR_79/S FILL
XFILL_1_OAI21X1_14 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_38_DFFSR_212 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_0_INVX1_155 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_0_DFFSR_70 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_0_INVX1_17 AND2X2_38/B DFFSR_59/S FILL
XFILL_17_DFFSR_63 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_28_DFFSR_23 AND2X2_38/B DFFSR_23/S FILL
XFILL_3_AND2X2_22 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_14_DFFSR_111 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_4_BUFX2_98 BUFX2_79/A DFFSR_7/S FILL
XFILL_7_NAND3X1_88 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_28_DFFSR_215 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_0_OAI21X1_17 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_11_OAI22X1_4 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_6_NAND3X1_91 AND2X2_38/B DFFSR_59/S FILL
XFILL_18_DFFSR_218 BUFX2_98/A DFFSR_32/S FILL
XFILL_5_NAND3X1_94 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_0_NAND3X1_137 BUFX2_7/gnd DFFSR_216/S FILL
XNAND3X1_91 BUFX2_93/A AND2X2_16/Y BUFX2_32/Y AND2X2_38/B AND2X2_22/A DFFSR_59/S NAND3X1
XFILL_4_NAND3X1_97 AND2X2_38/B DFFSR_59/S FILL
XFILL_33_DFFSR_2 BUFX2_79/A DFFSR_7/S FILL
XFILL_5_DFFPOSX1_11 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_0_DFFSR_108 OR2X2_6/gnd DFFSR_92/S FILL
XDFFSR_218 DFFSR_218/Q DFFSR_3/CLK BUFX2_65/Y DFFSR_32/S INVX1_71/A BUFX2_98/A DFFSR_32/S
+ DFFSR
XFILL_2_NAND2X1_173 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_41_DFFSR_139 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_25_DFFSR_70 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_36_DFFSR_30 BUFX2_98/A DFFSR_32/S FILL
XFILL_8_DFFSR_77 BUFX2_98/A DFFSR_32/S FILL
XFILL_4_DFFSR_215 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_31_DFFSR_142 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_45_DFFSR_246 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_21_DFFSR_145 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_35_DFFSR_249 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_14_DFFPOSX1_30 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_11_DFFSR_148 INVX1_67/gnd DFFSR_175/S FILL
XFILL_3_NAND2X1_107 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_25_DFFSR_252 AND2X2_38/B DFFSR_23/S FILL
XFILL_6_NOR2X1_24 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_15_DFFSR_255 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_0_NOR3X1_1 INVX1_3/gnd DFFSR_79/S FILL
XFILL_0_AOI22X1_10 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_10_OAI22X1_28 INVX1_3/gnd DFFSR_23/S FILL
XFILL_44_DFFSR_37 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_7_DFFSR_142 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_33_DFFSR_77 BUFX2_98/A DFFSR_32/S FILL
XFILL_24_DFFPOSX1_19 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_27_3_0 INVX1_3/gnd DFFSR_79/S FILL
XFILL_48_DFFSR_173 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_8_NAND3X1_49 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_9_OAI22X1_31 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_38_DFFSR_176 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_0_DFFSR_34 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_8_NAND3X1_222 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_0_INVX1_119 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_17_DFFSR_27 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_7_NAND3X1_52 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_1_DFFSR_252 AND2X2_38/B DFFSR_23/S FILL
XFILL_25_5_1 AND2X2_38/B DFFSR_23/S FILL
XFILL_8_OAI22X1_34 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_4_BUFX2_62 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_4_DFFPOSX1_41 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_28_DFFSR_179 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_6_NAND3X1_55 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_7_OAI22X1_37 INVX1_3/gnd DFFSR_23/S FILL
XFILL_7_4_0 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_18_DFFSR_182 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_5_NAND3X1_58 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_6_OAI22X1_40 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_0_NAND3X1_101 XOR2X1_4/gnd DFFSR_91/S FILL
XNAND3X1_55 NAND3X1_53/Y NAND3X1_55/B AOI22X1_7/Y OR2X2_3/gnd NOR2X1_26/B DFFSR_60/S
+ NAND3X1
XFILL_4_NAND3X1_61 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_41_DFFSR_84 BUFX2_99/A DFFSR_7/S FILL
XFILL_5_OAI22X1_43 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_5_6_1 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_3_NOR2X1_61 BUFX2_8/gnd DFFSR_51/S FILL
XOAI22X1_40 INVX1_97/Y OAI22X1_43/B INVX1_98/Y OAI22X1_43/D DFFSR_46/gnd NOR2X1_50/B
+ DFFSR_62/S OAI22X1
XFILL_5_OAI21X1_9 INVX1_67/gnd DFFSR_201/S FILL
XFILL_3_NAND3X1_64 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_4_OAI22X1_46 OR2X2_1/gnd DFFSR_59/S FILL
XDFFSR_182 INVX1_97/A CLKBUF1_31/Y BUFX2_60/Y DFFSR_208/S INVX1_98/A XOR2X1_1/gnd
+ DFFSR_208/S DFFSR
XFILL_2_NAND2X1_137 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_2_NAND3X1_67 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_41_DFFSR_103 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_3_OAI22X1_49 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_8_DFFSR_41 BUFX2_98/A DFFSR_6/S FILL
XFILL_25_DFFSR_34 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_14_DFFSR_74 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_4_DFFSR_179 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_1_NAND3X1_70 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_2_OAI22X1_52 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_31_DFFSR_106 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_45_DFFSR_210 BUFX2_98/A DFFSR_6/S FILL
XNAND2X1_3 NOR2X1_2/Y AND2X2_2/Y BUFX2_99/A OAI22X1_2/D DFFSR_7/S NAND2X1
XFILL_21_DFFSR_109 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_0_NAND3X1_73 INVX1_1/gnd DFFSR_97/S FILL
XFILL_35_DFFSR_213 INVX1_3/gnd DFFSR_23/S FILL
XFILL_0_OAI21X1_119 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_0_AND2X2_23 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_11_DFFSR_112 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_23_DFFPOSX1_49 BUFX2_99/A DFFSR_92/S FILL
XFILL_25_DFFSR_216 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_0_DFFSR_5 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_49_DFFSR_91 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_15_DFFSR_219 INVX1_67/gnd DFFSR_175/S FILL
XOAI22X1_2 INVX1_5/Y OAI22X1_2/B INVX1_6/Y OAI22X1_2/D NOR3X1_6/gnd NOR2X1_3/A DFFSR_79/S
+ OAI22X1
XINVX1_75 INVX1_75/A BUFX2_98/A INVX1_75/Y DFFSR_6/S INVX1
XFILL_5_DFFSR_88 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_33_DFFSR_41 BUFX2_98/A DFFSR_6/S FILL
XFILL_7_DFFSR_106 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_22_DFFSR_81 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_48_DFFSR_137 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_35_0_1 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_8_NAND3X1_13 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_8_NAND3X1_186 BUFX2_7/gnd DFFSR_151/S FILL
XINVX1_193 INVX1_193/A BUFX2_8/gnd INVX1_193/Y DFFSR_51/S INVX1
XFILL_38_DFFSR_140 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_18_5 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_1_DFFSR_216 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_7_NAND3X1_16 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_4_BUFX2_26 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_28_DFFSR_143 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_42_DFFSR_247 BUFX2_99/A DFFSR_7/S FILL
XFILL_33_2_2 INVX1_1/gnd DFFSR_53/S FILL
XFILL_1_NAND2X1_167 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_6_NAND3X1_19 BUFX2_99/A DFFSR_92/S FILL
XFILL_18_DFFSR_146 BUFX2_79/A DFFSR_7/S FILL
XFILL_32_DFFSR_250 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_14_NOR3X1_5 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_24_DFFSR_9 BUFX2_79/A DFFSR_6/S FILL
XFILL_5_NAND3X1_22 OR2X2_6/gnd DFFSR_53/S FILL
XNAND3X1_19 BUFX2_84/A AND2X2_3/Y BUFX2_20/Y BUFX2_99/A AND2X2_8/A DFFSR_92/S NAND3X1
XFILL_4_NAND3X1_25 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_22_DFFSR_253 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_2_INVX1_82 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_41_DFFSR_48 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_30_DFFSR_88 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_3_NOR2X1_25 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_13_DFFPOSX1_24 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_12_DFFSR_256 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_3_NAND3X1_28 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_4_OAI22X1_10 DFFSR_8/gnd DFFSR_60/S FILL
XDFFSR_146 INVX1_73/A CLKBUF1_3/Y BUFX2_65/Y DFFSR_7/S INVX1_74/A BUFX2_79/A DFFSR_7/S
+ DFFSR
XFILL_2_NAND2X1_101 INVX1_39/gnd DFFSR_54/S FILL
XFILL_2_NAND3X1_31 BUFX2_79/A DFFSR_6/S FILL
XFILL_3_OAI22X1_13 INVX1_1/gnd DFFSR_53/S FILL
XFILL_4_DFFSR_143 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_14_DFFSR_38 BUFX2_98/A DFFSR_6/S FILL
XFILL_1_NAND3X1_34 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_1_BUFX2_73 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_2_OAI22X1_16 AND2X2_38/B DFFSR_59/S FILL
XFILL_45_DFFSR_174 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_0_NAND3X1_37 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_8_DFFSR_250 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_1_OAI22X1_19 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_35_DFFSR_177 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_23_DFFPOSX1_13 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_0_OAI22X1_22 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_45_DFFSR_5 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_25_DFFSR_180 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_49_DFFSR_55 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_38_DFFSR_95 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_15_DFFSR_183 INVX1_67/gnd DFFSR_175/S FILL
XFILL_7_NAND3X1_216 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_3_DFFPOSX1_35 INVX1_39/gnd DFFSR_54/S FILL
XFILL_5_DFFSR_52 OR2X2_3/gnd DFFSR_4/S FILL
XDFFSR_92 DFFSR_92/Q DFFSR_92/CLK DFFSR_7/R DFFSR_92/S INVX1_26/A BUFX2_99/A DFFSR_92/S
+ DFFSR
XINVX1_39 DFFSR_62/Q INVX1_39/gnd INVX1_39/Y DFFSR_34/S INVX1
XFILL_11_DFFSR_85 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_22_DFFSR_45 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_0_NOR2X1_62 INVX1_67/gnd DFFSR_201/S FILL
XFILL_48_DFFSR_101 OR2X2_3/gnd DFFSR_4/S FILL
XINVX1_157 INVX1_157/A BUFX2_7/gnd INVX1_157/Y DFFSR_216/S INVX1
XFILL_38_DFFSR_104 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_8_NAND3X1_150 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_0_INVX1_7 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_1_DFFSR_180 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_28_DFFSR_107 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_42_DFFSR_211 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_1_NAND2X1_131 INVX1_3/gnd DFFSR_79/S FILL
XFILL_4_INVX1_154 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_7_AND2X2_21 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_18_DFFSR_110 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_32_DFFSR_214 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_1_NAND2X1_1 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_22_DFFSR_217 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_41_DFFSR_12 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_30_DFFSR_52 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_2_INVX1_46 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_2_DFFSR_99 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_19_DFFSR_92 BUFX2_99/A DFFSR_92/S FILL
XFILL_12_DFFSR_220 BUFX2_7/gnd DFFSR_151/S FILL
XDFFSR_110 DFFSR_118/D DFFSR_45/CLK DFFSR_35/R DFFSR_4/S DFFSR_110/D OR2X2_3/gnd DFFSR_4/S
+ DFFSR
XFILL_22_DFFPOSX1_43 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_4_DFFSR_107 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_6_NAND3X1_246 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_1_BUFX2_37 INVX1_1/gnd DFFSR_97/S FILL
XFILL_45_DFFSR_138 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_8_DFFSR_214 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_35_DFFSR_141 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_11_DFFSR_3 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_49_DFFSR_245 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_25_DFFSR_144 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_39_DFFSR_248 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_1_INVX1_191 INVX1_67/gnd DFFSR_175/S FILL
XFILL_49_DFFSR_19 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_27_DFFSR_99 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_38_DFFSR_59 AND2X2_38/B DFFSR_59/S FILL
XFILL_7_NAND3X1_180 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_15_DFFSR_147 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_29_DFFSR_251 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_0_NAND2X1_161 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_5_DFFSR_16 DFFSR_28/gnd DFFSR_3/S FILL
XDFFSR_56 DFFSR_16/D DFFSR_7/CLK DFFSR_9/R DFFSR_8/S DFFSR_56/D DFFSR_28/gnd DFFSR_8/S
+ DFFSR
XFILL_19_DFFSR_254 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_11_DFFSR_49 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_0_NOR2X1_26 DFFSR_8/gnd DFFSR_60/S FILL
XINVX1_121 INVX1_3/A DFFSR_34/gnd INVX1_121/Y DFFSR_1/S INVX1
XFILL_8_NAND3X1_114 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_12_DFFPOSX1_18 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_1_DFFSR_144 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_42_DFFSR_175 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_4_INVX1_118 BUFX2_98/A DFFSR_6/S FILL
XFILL_46_DFFSR_66 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_3_BUFX2_100 BUFX2_79/A DFFSR_6/S FILL
XFILL_5_DFFSR_251 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_32_DFFSR_178 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_22_DFFSR_181 INVX1_3/gnd DFFSR_79/S FILL
XFILL_30_DFFSR_16 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_2_DFFSR_63 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_2_INVX1_10 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_19_DFFSR_56 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_6_BUFX2_91 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_12_DFFSR_184 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_34_3_0 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_20_CLKBUF1_46 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_6_NAND3X1_210 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_45_DFFSR_102 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_32_5_1 INVX1_1/gnd DFFSR_97/S FILL
XFILL_2_DFFPOSX1_29 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_8_DFFSR_178 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_19_CLKBUF1_49 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_35_DFFSR_105 INVX1_1/gnd DFFSR_53/S FILL
XAND2X2_25 AND2X2_25/A AND2X2_25/B INVX1_39/gnd AND2X2_25/Y DFFSR_54/S AND2X2
XFILL_49_DFFSR_209 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_25_DFFSR_108 OR2X2_6/gnd DFFSR_92/S FILL
XNAND3X1_246 NAND2X1_113/Y NAND2X1_114/Y AOI21X1_43/Y OR2X2_4/gnd NAND3X1_246/Y DFFSR_3/S
+ NAND3X1
XFILL_39_DFFSR_212 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_1_INVX1_155 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_27_DFFSR_63 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_38_DFFSR_23 AND2X2_38/B DFFSR_23/S FILL
XFILL_4_AND2X2_22 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_15_DFFSR_111 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_7_NAND3X1_144 AND2X2_38/B DFFSR_59/S FILL
XFILL_29_DFFSR_215 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_11_DFFPOSX1_48 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_0_NAND2X1_125 OR2X2_2/gnd DFFSR_175/S FILL
XDFFSR_20 INVX1_28/A CLKBUF1_4/Y DFFSR_8/R DFFSR_5/S DFFSR_28/Q DFFSR_5/gnd DFFSR_5/S
+ DFFSR
XFILL_19_DFFSR_218 BUFX2_98/A DFFSR_32/S FILL
XFILL_11_DFFSR_13 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_1_DFFSR_108 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_21_DFFPOSX1_37 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_42_DFFSR_139 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_46_DFFSR_30 BUFX2_98/A DFFSR_32/S FILL
XFILL_35_DFFSR_70 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_5_DFFSR_215 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_32_DFFSR_142 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_5_NAND3X1_240 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_46_DFFSR_246 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_22_DFFSR_145 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_36_DFFSR_249 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_2_DFFSR_27 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_19_DFFSR_20 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_12_DFFSR_148 INVX1_67/gnd DFFSR_175/S FILL
XFILL_6_BUFX2_55 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_26_DFFSR_252 AND2X2_38/B DFFSR_23/S FILL
XFILL_42_0_1 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_16_DFFSR_255 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_1_NOR2X1_8 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_6_NAND3X1_174 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_8_DFFSR_142 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_19_CLKBUF1_13 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_43_DFFSR_77 BUFX2_98/A DFFSR_32/S FILL
XFILL_40_2_2 BUFX2_98/A DFFSR_6/S FILL
XFILL_18_CLKBUF1_16 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_49_DFFSR_173 XOR2X1_1/gnd DFFSR_208/S FILL
XNAND3X1_210 INVX1_164/A OAI21X1_69/Y OAI21X1_70/Y BUFX2_8/gnd NAND3X1_215/A DFFSR_81/S
+ NAND3X1
XFILL_39_DFFSR_176 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_17_CLKBUF1_19 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_1_INVX1_119 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_27_DFFSR_27 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_16_DFFSR_67 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_2_DFFSR_252 AND2X2_38/B DFFSR_23/S FILL
XFILL_7_NAND3X1_108 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_16_CLKBUF1_22 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_29_DFFSR_179 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_11_DFFPOSX1_12 AND2X2_38/B DFFSR_23/S FILL
XFILL_15_CLKBUF1_25 INVX1_67/gnd DFFSR_201/S FILL
XFILL_19_DFFSR_182 XOR2X1_1/gnd DFFSR_208/S FILL
XNOR2X1_64 NOR2X1_64/A NOR2X1_64/B AND2X2_38/B NOR2X1_64/Y DFFSR_59/S NOR2X1
XFILL_14_CLKBUF1_28 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_3_XOR2X1_4 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_13_CLKBUF1_31 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_23_DFFSR_6 BUFX2_79/A DFFSR_6/S FILL
XFILL_4_NOR2X1_61 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_6_OAI21X1_9 INVX1_67/gnd DFFSR_201/S FILL
XFILL_12_CLKBUF1_34 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_42_DFFSR_103 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_7_DFFSR_81 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_35_DFFSR_34 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_11_CLKBUF1_37 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_24_DFFSR_74 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_5_DFFSR_179 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_32_DFFSR_106 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_46_DFFSR_210 BUFX2_98/A DFFSR_6/S FILL
XFILL_10_CLKBUF1_40 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_5_NAND3X1_204 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_22_DFFSR_109 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_1_DFFPOSX1_23 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_36_DFFSR_213 INVX1_3/gnd DFFSR_23/S FILL
XFILL_1_AND2X2_23 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_6_BUFX2_19 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_12_DFFSR_112 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_26_DFFSR_216 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_9_CLKBUF1_43 AND2X2_38/B DFFSR_23/S FILL
XFILL_16_DFFSR_219 INVX1_67/gnd DFFSR_175/S FILL
XFILL_8_CLKBUF1_46 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_44_DFFSR_2 BUFX2_79/A DFFSR_7/S FILL
XFILL_6_NAND3X1_138 INVX1_67/gnd DFFSR_201/S FILL
XFILL_7_CLKBUF1_49 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_10_DFFPOSX1_42 INVX1_39/gnd DFFSR_34/S FILL
XFILL_43_DFFSR_41 BUFX2_98/A DFFSR_6/S FILL
XFILL_4_INVX1_75 BUFX2_98/A DFFSR_6/S FILL
XFILL_8_DFFSR_106 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_32_DFFSR_81 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_49_DFFSR_137 BUFX2_7/gnd DFFSR_216/S FILL
XNAND3X1_174 BUFX2_56/Y AND2X2_37/B NOR2X1_70/A NOR3X1_6/gnd NAND3X1_176/B DFFSR_79/S
+ NAND3X1
XFILL_39_DFFSR_140 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_16_DFFSR_31 BUFX2_79/A DFFSR_6/S FILL
XFILL_22_2 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_2_DFFSR_216 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_29_DFFSR_143 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_3_BUFX2_66 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_43_DFFSR_247 BUFX2_99/A DFFSR_7/S FILL
XFILL_20_DFFPOSX1_31 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_19_DFFSR_146 BUFX2_79/A DFFSR_7/S FILL
XFILL_33_DFFSR_250 DFFSR_8/gnd DFFSR_8/S FILL
XNOR2X1_28 NOR2X1_28/A OAI21X1_8/Y BUFX2_98/A NOR2X1_28/Y DFFSR_6/S NOR2X1
XFILL_4_NAND3X1_234 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_23_DFFSR_253 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_51_DFFSR_48 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_4_NOR2X1_25 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_40_DFFSR_88 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_13_DFFSR_256 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_7_DFFSR_45 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_13_DFFSR_78 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_24_DFFSR_38 BUFX2_98/A DFFSR_6/S FILL
XFILL_5_DFFSR_143 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_46_DFFSR_174 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_14_0_2 INVX1_39/gnd DFFSR_54/S FILL
XFILL_5_NAND3X1_168 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_9_DFFSR_250 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_36_DFFSR_177 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_26_DFFSR_180 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_48_DFFSR_95 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_8_CLKBUF1_10 INVX1_67/gnd DFFSR_201/S FILL
XFILL_16_DFFSR_183 INVX1_67/gnd DFFSR_175/S FILL
XFILL_6_NAND3X1_102 INVX1_3/gnd DFFSR_23/S FILL
XFILL_7_CLKBUF1_13 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_32_DFFSR_45 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_4_DFFSR_92 BUFX2_99/A DFFSR_92/S FILL
XFILL_21_DFFSR_85 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_1_NOR2X1_62 INVX1_67/gnd DFFSR_201/S FILL
XFILL_6_CLKBUF1_16 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_49_DFFSR_101 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_5_CLKBUF1_19 BUFX2_8/gnd DFFSR_81/S FILL
XNAND3X1_138 INVX1_131/Y OAI21X1_26/C OR2X2_2/Y INVX1_67/gnd OAI21X1_23/C DFFSR_201/S
+ NAND3X1
XFILL_39_DFFSR_104 DFFSR_28/gnd DFFSR_8/S FILL
XCLKBUF1_16 BUFX2_2/Y OR2X2_3/gnd DFFSR_57/CLK DFFSR_4/S CLKBUF1
XFILL_5_6 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_4_CLKBUF1_22 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_3_BUFX2_30 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_2_DFFSR_180 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_29_DFFSR_107 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_43_DFFSR_211 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_3_CLKBUF1_25 INVX1_67/gnd DFFSR_201/S FILL
XFILL_8_AND2X2_21 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_19_DFFSR_110 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_41_3_0 BUFX2_98/A DFFSR_32/S FILL
XFILL_33_DFFSR_214 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_2_CLKBUF1_28 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_2_NAND2X1_1 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_23_DFFSR_217 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_1_CLKBUF1_31 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_4_NAND3X1_198 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_40_DFFSR_52 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_39_5_1 BUFX2_79/A DFFSR_6/S FILL
XFILL_29_DFFSR_92 BUFX2_99/A DFFSR_92/S FILL
XFILL_1_INVX1_86 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_0_CLKBUF1_34 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_13_DFFSR_220 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_0_DFFPOSX1_17 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_13_DFFSR_42 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_5_DFFSR_107 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_0_BUFX2_77 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_5_NAND3X1_132 AND2X2_38/B DFFSR_23/S FILL
XFILL_46_DFFSR_138 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_9_DFFSR_214 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_36_DFFSR_141 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_50_DFFSR_245 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_35_DFFSR_9 BUFX2_79/A DFFSR_6/S FILL
XFILL_26_DFFSR_144 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_40_DFFSR_248 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_2_INVX1_191 INVX1_67/gnd DFFSR_175/S FILL
XFILL_37_DFFSR_99 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_48_DFFSR_59 AND2X2_38/B DFFSR_59/S FILL
XFILL_44_2 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_16_DFFSR_147 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_30_DFFSR_251 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_20_DFFSR_254 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_4_DFFSR_56 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_21_DFFSR_49 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_19_DFFPOSX1_25 BUFX2_79/A DFFSR_6/S FILL
XFILL_10_DFFSR_89 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_1_NOR2X1_26 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_10_DFFSR_257 INVX1_39/gnd DFFSR_34/S FILL
XNAND3X1_102 DFFSR_205/D BUFX2_29/Y NOR2X1_31/Y INVX1_3/gnd NAND3X1_103/B DFFSR_23/S
+ NAND3X1
XFILL_3_NAND3X1_228 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_2_DFFSR_144 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_43_DFFSR_175 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_4_BUFX2_100 BUFX2_79/A DFFSR_6/S FILL
XFILL_6_DFFSR_251 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_33_DFFSR_178 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_49_0_1 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_23_DFFSR_181 INVX1_3/gnd DFFSR_79/S FILL
XFILL_4_NAND3X1_162 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_1_INVX1_50 BUFX2_98/A DFFSR_6/S FILL
XFILL_40_DFFSR_16 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_29_DFFSR_56 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_18_DFFSR_96 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_13_DFFSR_184 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_47_2_2 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_9_DFFPOSX1_36 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_0_BUFX2_41 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_46_DFFSR_102 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_9_DFFSR_178 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_36_DFFSR_105 INVX1_1/gnd DFFSR_53/S FILL
XFILL_50_DFFSR_209 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_26_DFFSR_108 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_40_DFFSR_212 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_2_INVX1_155 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_37_DFFSR_63 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_48_DFFSR_23 AND2X2_38/B DFFSR_23/S FILL
XFILL_5_AND2X2_22 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_16_DFFSR_111 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_30_DFFSR_215 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_15_1_0 INVX1_39/gnd DFFSR_34/S FILL
XFILL_20_DFFSR_218 BUFX2_98/A DFFSR_32/S FILL
XFILL_4_DFFSR_20 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_21_DFFSR_13 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_10_DFFSR_53 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_5_OAI21X1_114 AND2X2_38/B DFFSR_59/S FILL
XFILL_10_DFFSR_221 AND2X2_38/B DFFSR_59/S FILL
XFILL_13_3_1 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_3_NAND3X1_192 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_3_NOR2X1_1 BUFX2_99/A DFFSR_92/S FILL
XFILL_2_DFFSR_108 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_11_5_2 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_22_DFFSR_3 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_43_DFFSR_139 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_45_DFFSR_70 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_6_DFFSR_215 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_33_DFFSR_142 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_47_DFFSR_246 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_23_DFFSR_145 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_4_NAND3X1_126 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_37_DFFSR_249 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_1_INVX1_14 BUFX2_98/A DFFSR_6/S FILL
XFILL_18_DFFSR_60 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_29_DFFSR_20 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_1_DFFSR_67 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_13_DFFSR_148 INVX1_67/gnd DFFSR_175/S FILL
XFILL_5_BUFX2_95 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_6_BUFX2_4 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_27_DFFSR_252 AND2X2_38/B DFFSR_23/S FILL
XFILL_6_NAND2X1_162 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_49_7 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_17_DFFSR_255 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_9_DFFSR_142 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_18_DFFPOSX1_19 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_50_DFFSR_173 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_19_DFFPOSX1_1 INVX1_39/gnd DFFSR_34/S FILL
XFILL_40_DFFSR_176 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_37_DFFSR_27 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_9_DFFSR_74 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_2_INVX1_119 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_26_DFFSR_67 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_2_NAND3X1_222 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_3_DFFSR_252 AND2X2_38/B DFFSR_23/S FILL
XFILL_18_DFFPOSX1_4 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_30_DFFSR_179 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_17_DFFPOSX1_7 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_20_DFFSR_182 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_10_DFFSR_17 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_10_DFFSR_185 INVX1_39/gnd DFFSR_54/S FILL
XFILL_21_0_2 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_3_NAND3X1_156 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_5_NOR2X1_61 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_7_OAI21X1_9 INVX1_67/gnd DFFSR_201/S FILL
XFILL_43_DFFSR_103 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_8_DFFPOSX1_30 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_34_DFFSR_74 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_45_DFFSR_34 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_6_DFFSR_179 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_33_DFFSR_106 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_47_DFFSR_210 BUFX2_98/A DFFSR_6/S FILL
XFILL_1_1_2 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_23_DFFSR_109 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_37_DFFSR_213 INVX1_3/gnd DFFSR_23/S FILL
XFILL_18_DFFSR_24 BUFX2_98/A DFFSR_6/S FILL
XFILL_1_DFFSR_31 BUFX2_79/A DFFSR_6/S FILL
XFILL_2_AND2X2_23 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_13_DFFSR_112 OR2X2_4/gnd DFFSR_32/S FILL
XBUFX2_99 BUFX2_99/A BUFX2_99/A BUFX2_99/Y DFFSR_7/S BUFX2
XFILL_5_BUFX2_59 AND2X2_38/B DFFSR_23/S FILL
XFILL_17_DFFPOSX1_49 BUFX2_99/A DFFSR_92/S FILL
XFILL_27_DFFSR_216 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_10_OAI22X1_5 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_6_NAND2X1_126 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_17_DFFSR_219 INVX1_67/gnd DFFSR_175/S FILL
XFILL_9_NOR3X1_5 BUFX2_7/gnd DFFSR_216/S FILL
XXOR2X1_1 XOR2X1_1/A XOR2X1_1/B XOR2X1_1/gnd XOR2X1_1/Y DFFSR_208/S XOR2X1
XFILL_42_DFFSR_81 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_9_DFFSR_106 XOR2X1_4/gnd DFFSR_91/S FILL
XNAND2X1_162 DFFPOSX1_29/Q INVX1_208/Y BUFX2_72/gnd AOI21X1_57/A DFFSR_201/S NAND2X1
XFILL_48_3_0 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_50_DFFSR_137 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_4_OAI21X1_108 INVX1_1/gnd DFFSR_53/S FILL
XFILL_8_AOI21X1_54 AND2X2_38/B DFFSR_59/S FILL
XFILL_27_DFFPOSX1_38 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_40_DFFSR_140 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_7_AOI21X1_57 INVX1_67/gnd DFFSR_201/S FILL
XFILL_9_DFFSR_38 BUFX2_98/A DFFSR_6/S FILL
XFILL_26_DFFSR_31 BUFX2_79/A DFFSR_6/S FILL
XFILL_2_NAND3X1_186 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_15_DFFSR_71 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_3_DFFSR_216 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_30_DFFSR_143 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_46_5_1 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_6_AOI21X1_60 BUFX2_79/A DFFSR_7/S FILL
XFILL_44_DFFSR_247 BUFX2_99/A DFFSR_7/S FILL
XFILL_20_DFFSR_146 BUFX2_79/A DFFSR_7/S FILL
XFILL_5_AOI21X1_63 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_34_DFFSR_250 DFFSR_8/gnd DFFSR_8/S FILL
XAOI21X1_60 AOI21X1_60/A AOI21X1_60/B BUFX2_40/Y BUFX2_79/A AOI21X1_60/Y DFFSR_7/S
+ AOI21X1
XFILL_10_DFFSR_149 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_2_XOR2X1_8 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_4_AOI21X1_66 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_24_DFFSR_253 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_50_DFFSR_88 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_5_NOR2X1_25 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_3_AOI21X1_69 INVX1_1/gnd DFFSR_97/S FILL
XFILL_3_NAND3X1_120 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_14_DFFSR_256 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_5_NAND2X1_156 AND2X2_38/B DFFSR_59/S FILL
XFILL_6_DFFSR_85 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_23_DFFSR_78 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_34_DFFSR_38 BUFX2_98/A DFFSR_6/S FILL
XFILL_6_DFFSR_143 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_47_DFFSR_174 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_37_DFFSR_177 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_8_OR2X2_2 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_5_BUFX2_23 XOR2X1_1/gnd DFFSR_151/S FILL
XBUFX2_63 BUFX2_60/A BUFX2_98/A BUFX2_63/Y DFFSR_32/S BUFX2
XFILL_0_DFFSR_253 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_17_DFFPOSX1_13 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_12_6_0 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_27_DFFSR_180 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_9_OAI21X1_99 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_17_DFFSR_183 INVX1_67/gnd DFFSR_175/S FILL
XFILL_34_DFFSR_6 BUFX2_79/A DFFSR_6/S FILL
XFILL_15_NOR3X1_2 INVX1_1/gnd DFFSR_53/S FILL
XFILL_1_NAND3X1_216 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_42_DFFSR_45 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_3_INVX1_79 INVX1_39/gnd DFFSR_54/S FILL
XFILL_31_DFFSR_85 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_9_AOI21X1_15 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_2_NOR2X1_62 INVX1_67/gnd DFFSR_201/S FILL
XNAND2X1_126 BUFX2_53/Y AOI21X1_7/C OR2X2_2/gnd OAI21X1_95/C DFFSR_175/S NAND2X1
XFILL_50_DFFSR_101 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_8_AOI21X1_18 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_7_DFFPOSX1_1 INVX1_39/gnd DFFSR_34/S FILL
XFILL_40_DFFSR_104 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_9_3 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_7_AOI21X1_21 INVX1_39/gnd DFFSR_54/S FILL
XFILL_6_DFFPOSX1_4 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_15_DFFSR_35 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_2_NAND3X1_150 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_3_DFFSR_180 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_2_BUFX2_70 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_30_DFFSR_107 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_5_DFFPOSX1_7 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_44_DFFSR_211 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_6_AOI21X1_24 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_54_2_2 DFFSR_5/gnd DFFSR_5/S FILL
XDFFPOSX1_4 INVX1_120/A CLKBUF1_44/Y AND2X2_27/Y DFFSR_62/gnd DFFSR_62/S DFFPOSX1
XFILL_20_DFFSR_110 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_7_DFFPOSX1_24 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_5_AOI21X1_27 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_34_DFFSR_214 BUFX2_72/gnd DFFSR_276/S FILL
XAOI21X1_24 NAND2X1_90/A NAND2X1_90/B INVX1_162/A DFFSR_46/gnd OAI21X1_74/A DFFSR_54/S
+ AOI21X1
XFILL_10_DFFSR_113 BUFX2_99/A DFFSR_92/S FILL
XFILL_3_NAND2X1_1 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_4_AOI21X1_30 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_24_DFFSR_217 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_50_DFFSR_52 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_39_DFFSR_92 BUFX2_99/A DFFSR_92/S FILL
XFILL_3_AOI21X1_33 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_14_DFFSR_220 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_16_DFFPOSX1_43 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_2_AOI21X1_36 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_0_AND2X2_1 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_5_NAND2X1_120 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_23_DFFSR_42 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_6_DFFSR_49 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_1_AOI21X1_39 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_12_DFFSR_82 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_6_DFFSR_107 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_0_NAND3X1_246 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_47_DFFSR_138 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_0_AOI21X1_42 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_22_1_0 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_37_DFFSR_141 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_51_DFFSR_245 DFFSR_34/gnd DFFSR_34/S FILL
XBUFX2_27 BUFX2_27/A DFFSR_62/gnd BUFX2_27/Y DFFSR_208/S BUFX2
XFILL_0_DFFSR_217 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_3_OAI21X1_102 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_27_DFFSR_144 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_26_DFFPOSX1_32 INVX1_67/gnd DFFSR_201/S FILL
XFILL_41_DFFSR_248 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_9_OAI21X1_63 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_31_4 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_3_INVX1_191 INVX1_67/gnd DFFSR_175/S FILL
XFILL_47_DFFSR_99 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_20_3_1 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_17_DFFSR_147 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_8_OAI21X1_66 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_31_DFFSR_251 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_1_NAND3X1_180 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_2_2_0 INVX1_67/gnd DFFSR_201/S FILL
XFILL_6_NAND2X1_87 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_7_OAI21X1_69 INVX1_3/gnd DFFSR_23/S FILL
XFILL_8_AND2X2_8 BUFX2_99/A DFFSR_7/S FILL
XFILL_21_DFFSR_254 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_3_INVX1_43 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_3_DFFSR_96 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_18_5_2 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_31_DFFSR_49 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_20_DFFSR_89 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_2_NOR2X1_26 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_6_OAI21X1_72 INVX1_3/gnd DFFSR_23/S FILL
XFILL_11_DFFSR_257 INVX1_39/gnd DFFSR_34/S FILL
XFILL_5_NAND2X1_90 DFFSR_46/gnd DFFSR_54/S FILL
XNAND2X1_87 BUFX2_57/Y AND2X2_37/B NOR3X1_6/gnd NOR2X1_70/B DFFSR_91/S NAND2X1
XFILL_0_4_1 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_4_NAND2X1_93 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_5_OAI21X1_75 INVX1_39/gnd DFFSR_54/S FILL
XOAI21X1_72 OR2X2_3/A OAI21X1_72/B OAI21X1_61/Y INVX1_3/gnd OAI21X1_72/Y DFFSR_23/S
+ OAI21X1
XFILL_2_NAND3X1_114 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_4_OAI21X1_78 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_3_NAND2X1_96 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_3_DFFSR_144 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_2_BUFX2_34 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_44_DFFSR_175 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_2_NAND2X1_99 INVX1_39/gnd DFFSR_54/S FILL
XFILL_3_OAI21X1_81 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_5_BUFX2_100 BUFX2_79/A DFFSR_6/S FILL
XFILL_7_DFFSR_251 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_1_DFFSR_9 BUFX2_79/A DFFSR_6/S FILL
XFILL_34_DFFSR_178 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_4_NAND2X1_150 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_2_OAI21X1_84 BUFX2_98/A DFFSR_6/S FILL
XFILL_24_DFFSR_181 INVX1_3/gnd DFFSR_79/S FILL
XFILL_1_OAI21X1_87 BUFX2_79/A DFFSR_7/S FILL
XFILL_50_DFFSR_16 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_39_DFFSR_56 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_28_DFFSR_96 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_0_INVX1_90 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_14_DFFSR_184 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_0_OAI21X1_90 BUFX2_98/A DFFSR_32/S FILL
XFILL_6_DFFSR_13 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_12_DFFSR_46 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_5_BUFX2_1 OR2X2_4/gnd DFFSR_32/S FILL
XBUFX2_5 BUFX2_3/A AND2X2_38/B BUFX2_5/Y DFFSR_59/S BUFX2
XFILL_47_DFFSR_102 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_0_NAND3X1_210 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_37_DFFSR_105 INVX1_1/gnd DFFSR_53/S FILL
XFILL_0_DFFSR_181 INVX1_3/gnd DFFSR_79/S FILL
XFILL_27_DFFSR_108 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_41_DFFSR_212 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_3_INVX1_155 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_47_DFFSR_63 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_6_AND2X2_22 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_17_DFFSR_111 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_28_0_2 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_8_OAI21X1_30 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_1_NAND3X1_144 AND2X2_38/B DFFSR_59/S FILL
XFILL_31_DFFSR_215 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_0_NAND2X1_2 BUFX2_99/A DFFSR_7/S FILL
XFILL_6_NAND2X1_51 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_7_OAI21X1_33 INVX1_3/gnd DFFSR_79/S FILL
XFILL_21_DFFSR_218 BUFX2_98/A DFFSR_32/S FILL
XFILL_3_DFFSR_60 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_31_DFFSR_13 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_20_DFFSR_53 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_6_DFFPOSX1_18 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_3_NAND2X1_180 INVX1_1/gnd DFFSR_97/S FILL
XFILL_5_NAND2X1_54 AND2X2_38/B DFFSR_59/S FILL
XFILL_11_DFFSR_221 AND2X2_38/B DFFSR_59/S FILL
XFILL_6_OAI21X1_36 BUFX2_8/gnd DFFSR_51/S FILL
XNAND2X1_51 DFFSR_240/Q NOR2X1_34/Y XOR2X1_4/gnd OAI21X1_16/C DFFSR_97/S NAND2X1
XFILL_4_NAND2X1_57 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_5_OAI21X1_39 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_8_1_2 XOR2X1_1/gnd DFFSR_151/S FILL
XOAI21X1_36 INVX1_133/Y INVX1_150/Y OAI21X1_36/C BUFX2_8/gnd OAI21X1_37/C DFFSR_51/S
+ OAI21X1
XFILL_4_OAI21X1_42 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_3_DFFSR_108 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_3_NAND2X1_60 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_0_OAI22X1_1 INVX1_1/gnd DFFSR_53/S FILL
XFILL_44_DFFSR_139 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_2_NAND2X1_63 AND2X2_38/B DFFSR_59/S FILL
XFILL_15_DFFPOSX1_37 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_46_DFFSR_9 BUFX2_79/A DFFSR_6/S FILL
XFILL_3_OAI21X1_45 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_7_DFFSR_215 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_34_DFFSR_142 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_4_NAND2X1_114 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_2_OAI21X1_48 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_1_NAND2X1_66 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_48_DFFSR_246 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_11_AOI22X1_14 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_24_DFFSR_145 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_0_NAND2X1_69 INVX1_3/gnd DFFSR_23/S FILL
XFILL_1_OAI21X1_51 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_38_DFFSR_249 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_0_INVX1_192 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_28_DFFSR_60 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_0_INVX1_54 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_39_DFFSR_20 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_10_AOI22X1_17 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_14_DFFSR_148 INVX1_67/gnd DFFSR_175/S FILL
XFILL_0_OAI21X1_54 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_28_DFFSR_252 AND2X2_38/B DFFSR_23/S FILL
XFILL_53_4 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_18_DFFSR_255 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_25_DFFPOSX1_26 AND2X2_38/B DFFSR_23/S FILL
XFILL_12_DFFSR_10 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_9_AOI22X1_20 INVX1_39/gnd DFFSR_34/S FILL
XFILL_0_NAND3X1_174 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_8_AOI22X1_23 INVX1_39/gnd DFFSR_34/S FILL
XFILL_53_5_1 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_9_NAND3X1_229 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_7_AOI22X1_26 INVX1_1/gnd DFFSR_97/S FILL
XFILL_5_DFFPOSX1_48 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_51_DFFSR_173 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_0_DFFSR_145 BUFX2_72/gnd DFFSR_201/S FILL
XDFFSR_255 BUFX2_96/A DFFSR_3/CLK BUFX2_65/Y DFFSR_32/S INVX1_110/A OR2X2_4/gnd DFFSR_32/S
+ DFFSR
XFILL_6_AOI22X1_29 INVX1_1/gnd DFFSR_53/S FILL
XFILL_41_DFFSR_176 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_47_DFFSR_27 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_3_INVX1_119 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_36_DFFSR_67 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_4_DFFSR_252 AND2X2_38/B DFFSR_23/S FILL
XFILL_31_DFFSR_179 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_1_NAND3X1_108 BUFX2_8/gnd DFFSR_81/S FILL
XAOI22X1_29 AOI22X1_26/A AOI22X1_26/B AOI22X1_29/C INVX1_174/A INVX1_1/gnd OAI21X1_72/B
+ DFFSR_53/S AOI22X1
XFILL_6_NAND2X1_15 BUFX2_99/A DFFSR_92/S FILL
XFILL_21_DFFSR_182 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_3_DFFSR_24 BUFX2_98/A DFFSR_6/S FILL
XFILL_20_DFFSR_17 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_5_NAND2X1_18 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_11_DFFSR_185 INVX1_39/gnd DFFSR_54/S FILL
XFILL_3_NAND2X1_144 DFFSR_46/gnd DFFSR_62/S FILL
XNAND2X1_15 DFFSR_115/D NOR2X1_5/Y BUFX2_99/A OAI21X1_3/C DFFSR_92/S NAND2X1
XFILL_4_NAND2X1_21 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_6_NOR2X1_61 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_8_OAI21X1_9 INVX1_67/gnd DFFSR_201/S FILL
XFILL_3_NAND2X1_24 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_2_NOR2X1_5 OR2X2_6/gnd DFFSR_53/S FILL
XDFFPOSX1_18 INVX1_154/A CLKBUF1_49/Y OAI21X1_45/Y DFFSR_46/gnd DFFSR_62/S DFFPOSX1
XFILL_44_DFFSR_103 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_12_DFFSR_7 BUFX2_79/A DFFSR_7/S FILL
XFILL_2_NAND2X1_27 AND2X2_38/B DFFSR_23/S FILL
XFILL_19_6_0 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_44_DFFSR_74 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_7_DFFSR_179 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_34_DFFSR_106 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_48_DFFSR_210 BUFX2_98/A DFFSR_6/S FILL
XFILL_1_NAND2X1_30 AND2X2_38/B DFFSR_23/S FILL
XFILL_2_OAI21X1_12 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_24_DFFSR_109 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_8_NAND3X1_86 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_0_NAND2X1_33 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_1_OAI21X1_15 INVX1_3/gnd DFFSR_79/S FILL
XFILL_28_DFFSR_24 BUFX2_98/A DFFSR_6/S FILL
XFILL_0_DFFSR_71 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_38_DFFSR_213 INVX1_3/gnd DFFSR_23/S FILL
XFILL_0_INVX1_18 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_0_INVX1_156 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_17_DFFSR_64 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_3_AND2X2_23 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_14_DFFSR_112 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_7_NAND3X1_89 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_4_BUFX2_99 BUFX2_99/A DFFSR_7/S FILL
XFILL_0_OAI21X1_18 INVX1_39/gnd DFFSR_34/S FILL
XFILL_28_DFFSR_216 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_11_OAI22X1_5 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_6_NAND3X1_92 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_18_DFFSR_219 INVX1_67/gnd DFFSR_175/S FILL
XFILL_5_NAND3X1_95 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_0_NAND3X1_138 INVX1_67/gnd DFFSR_201/S FILL
XNAND3X1_92 NAND2X1_44/Y NAND3X1_89/Y AND2X2_22/Y DFFSR_34/gnd NOR2X1_46/A DFFSR_1/S
+ NAND3X1
XFILL_4_XOR2X1_1 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_4_NAND3X1_98 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_33_DFFSR_3 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_51_DFFSR_137 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_5_DFFPOSX1_12 AND2X2_38/B DFFSR_23/S FILL
XDFFSR_219 DFFSR_219/Q CLKBUF1_25/Y BUFX2_60/Y DFFSR_175/S INVX1_78/A INVX1_67/gnd
+ DFFSR_175/S DFFSR
XFILL_0_DFFSR_109 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_13_1 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_2_NAND2X1_174 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_41_DFFSR_140 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_8_DFFSR_78 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_36_DFFSR_31 BUFX2_79/A DFFSR_6/S FILL
XFILL_25_DFFSR_71 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_4_DFFSR_216 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_31_DFFSR_143 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_45_DFFSR_247 BUFX2_99/A DFFSR_7/S FILL
XFILL_21_DFFSR_146 BUFX2_79/A DFFSR_7/S FILL
XFILL_14_DFFPOSX1_31 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_35_DFFSR_250 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_11_DFFSR_149 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_3_NAND2X1_108 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_25_DFFSR_253 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_6_NOR2X1_25 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_15_DFFSR_256 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_29_1_0 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_0_NOR3X1_2 INVX1_1/gnd DFFSR_53/S FILL
XFILL_0_AOI22X1_11 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_10_OAI22X1_29 INVX1_3/gnd DFFSR_79/S FILL
XFILL_33_DFFSR_78 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_44_DFFSR_38 BUFX2_98/A DFFSR_6/S FILL
XFILL_7_DFFSR_143 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_27_3_1 INVX1_3/gnd DFFSR_79/S FILL
XFILL_24_DFFPOSX1_20 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_48_DFFSR_174 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_8_NAND3X1_50 BUFX2_98/A DFFSR_6/S FILL
XFILL_9_OAI22X1_32 INVX1_39/gnd DFFSR_54/S FILL
XFILL_38_DFFSR_177 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_9_2_0 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_0_DFFSR_35 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_8_NAND3X1_223 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_0_INVX1_120 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_17_DFFSR_28 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_7_NAND3X1_53 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_25_5_2 AND2X2_38/B DFFSR_23/S FILL
XFILL_8_OAI22X1_35 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_1_DFFSR_253 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_4_BUFX2_63 BUFX2_98/A DFFSR_32/S FILL
XFILL_28_DFFSR_180 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_4_DFFPOSX1_42 INVX1_39/gnd DFFSR_34/S FILL
XFILL_6_NAND3X1_56 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_7_OAI22X1_38 AND2X2_38/B DFFSR_23/S FILL
XFILL_18_DFFSR_183 INVX1_67/gnd DFFSR_175/S FILL
XFILL_7_4_1 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_5_NAND3X1_59 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_6_OAI22X1_41 INVX1_39/gnd DFFSR_54/S FILL
XNAND3X1_56 NOR2X1_24/Y NOR2X1_25/Y NOR2X1_26/Y DFFSR_28/gnd XOR2X1_15/A DFFSR_8/S
+ NAND3X1
XFILL_0_NAND3X1_102 INVX1_3/gnd DFFSR_23/S FILL
XFILL_4_NAND3X1_62 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_5_OAI22X1_44 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_41_DFFSR_85 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_3_NOR2X1_62 INVX1_67/gnd DFFSR_201/S FILL
XFILL_5_6_2 OR2X2_2/gnd DFFSR_216/S FILL
XOAI22X1_41 INVX1_99/Y OAI22X1_41/B INVX1_100/Y OAI22X1_41/D INVX1_39/gnd NOR2X1_50/A
+ DFFSR_54/S OAI22X1
XFILL_51_DFFSR_101 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_4_OAI22X1_47 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_3_NAND3X1_65 DFFSR_62/gnd DFFSR_208/S FILL
XDFFSR_183 DFFSR_183/Q CLKBUF1_34/Y BUFX2_62/Y DFFSR_175/S DFFSR_183/D INVX1_67/gnd
+ DFFSR_175/S DFFSR
XFILL_2_NAND2X1_138 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_41_DFFSR_104 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_2_NAND3X1_68 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_8_DFFSR_42 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_3_OAI22X1_50 INVX1_3/gnd DFFSR_23/S FILL
XFILL_25_DFFSR_35 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_14_DFFSR_75 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_4_DFFSR_180 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_1_NAND3X1_71 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_31_DFFSR_107 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_45_DFFSR_211 BUFX2_7/gnd DFFSR_216/S FILL
XNAND2X1_4 NOR2X1_1/Y NOR2X1_2/Y BUFX2_98/A OAI22X1_2/B DFFSR_6/S NAND2X1
XFILL_21_DFFSR_110 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_0_NAND3X1_74 INVX1_1/gnd DFFSR_97/S FILL
XFILL_35_DFFSR_214 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_23_DFFPOSX1_50 INVX1_1/gnd DFFSR_53/S FILL
XFILL_0_AND2X2_24 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_11_DFFSR_113 BUFX2_99/A DFFSR_92/S FILL
XFILL_4_NAND2X1_1 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_25_DFFSR_217 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_0_DFFSR_6 BUFX2_79/A DFFSR_6/S FILL
XFILL_49_DFFSR_92 BUFX2_99/A DFFSR_92/S FILL
XFILL_15_DFFSR_220 BUFX2_7/gnd DFFSR_151/S FILL
XOAI22X1_3 INVX1_7/Y OAI22X1_6/B INVX1_8/Y OAI22X1_6/D OR2X2_4/gnd NOR2X1_6/A DFFSR_3/S
+ OAI22X1
XINVX1_76 INVX1_76/A DFFSR_1/gnd INVX1_76/Y DFFSR_1/S INVX1
XFILL_33_DFFSR_42 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_5_DFFSR_89 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_22_DFFSR_82 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_7_DFFSR_107 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_9_NAND3X1_11 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_48_DFFSR_138 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_35_0_2 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_8_NAND3X1_14 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_38_DFFSR_141 XOR2X1_4/gnd DFFSR_91/S FILL
XINVX1_194 INVX1_194/A BUFX2_72/gnd INVX1_194/Y DFFSR_276/S INVX1
XFILL_8_NAND3X1_187 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_1_DFFSR_217 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_7_NAND3X1_17 BUFX2_99/A DFFSR_7/S FILL
XFILL_18_6 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_4_BUFX2_27 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_35_1 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_28_DFFSR_144 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_1_NAND2X1_168 BUFX2_79/A DFFSR_6/S FILL
XFILL_42_DFFSR_248 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_6_NAND3X1_20 BUFX2_99/A DFFSR_7/S FILL
XFILL_18_DFFSR_147 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_32_DFFSR_251 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_14_NOR3X1_6 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_5_NAND3X1_23 OR2X2_6/gnd DFFSR_53/S FILL
XNAND3X1_20 NAND3X1_20/A NAND3X1_17/Y AND2X2_8/Y BUFX2_99/A NOR2X1_14/A DFFSR_7/S
+ NAND3X1
XFILL_22_DFFSR_254 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_4_NAND3X1_26 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_9_NAND3X1_121 INVX1_1/gnd DFFSR_97/S FILL
XFILL_41_DFFSR_49 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_30_DFFSR_89 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_2_INVX1_83 INVX1_39/gnd DFFSR_54/S FILL
XFILL_3_NOR2X1_26 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_13_DFFPOSX1_25 BUFX2_79/A DFFSR_6/S FILL
XFILL_12_DFFSR_257 INVX1_39/gnd DFFSR_34/S FILL
XFILL_3_NAND3X1_29 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_4_OAI22X1_11 BUFX2_99/A DFFSR_92/S FILL
XFILL_2_NAND2X1_102 OR2X2_1/gnd DFFSR_51/S FILL
XDFFSR_147 INVX1_80/A CLKBUF1_17/Y BUFX2_69/Y DFFSR_1/S INVX1_81/A DFFSR_1/gnd DFFSR_1/S
+ DFFSR
XFILL_3_OAI22X1_14 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_2_NAND3X1_32 BUFX2_79/A DFFSR_7/S FILL
XFILL_14_DFFSR_39 INVX1_3/gnd DFFSR_79/S FILL
XFILL_4_DFFSR_144 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_1_BUFX2_74 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_1_NAND3X1_35 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_2_OAI22X1_17 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_45_DFFSR_175 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_6_BUFX2_100 BUFX2_79/A DFFSR_6/S FILL
XFILL_8_DFFSR_251 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_1_OAI22X1_20 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_0_NAND3X1_38 BUFX2_98/A DFFSR_32/S FILL
XFILL_35_DFFSR_178 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_23_DFFPOSX1_14 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_0_OAI22X1_23 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_45_DFFSR_6 BUFX2_79/A DFFSR_6/S FILL
XFILL_25_DFFSR_181 INVX1_3/gnd DFFSR_79/S FILL
XFILL_49_DFFSR_56 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_38_DFFSR_96 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_15_DFFSR_184 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_7_NAND3X1_217 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_3_DFFPOSX1_36 OR2X2_2/gnd DFFSR_175/S FILL
XDFFSR_93 DFFSR_93/Q DFFSR_93/CLK DFFSR_5/R DFFSR_60/S INVX1_33/A OR2X2_3/gnd DFFSR_60/S
+ DFFSR
XINVX1_40 DFFSR_86/Q DFFSR_4/gnd INVX1_40/Y DFFSR_98/S INVX1
XFILL_5_DFFSR_53 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_11_DFFSR_86 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_22_DFFSR_46 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_0_NOR2X1_63 INVX1_3/gnd DFFSR_23/S FILL
XFILL_48_DFFSR_102 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_38_DFFSR_105 INVX1_1/gnd DFFSR_53/S FILL
XFILL_8_NAND3X1_151 DFFSR_1/gnd DFFSR_81/S FILL
XINVX1_158 INVX1_158/A INVX1_39/gnd INVX1_158/Y DFFSR_34/S INVX1
XFILL_0_INVX1_8 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_1_DFFSR_181 INVX1_3/gnd DFFSR_79/S FILL
XFILL_28_DFFSR_108 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_1_NAND2X1_132 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_42_DFFSR_212 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_4_INVX1_155 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_7_AND2X2_22 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_18_DFFSR_111 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_32_DFFSR_215 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_1_NAND2X1_2 BUFX2_99/A DFFSR_7/S FILL
XFILL_22_DFFSR_218 BUFX2_98/A DFFSR_32/S FILL
XFILL_19_DFFSR_93 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_2_INVX1_47 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_41_DFFSR_13 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_30_DFFSR_53 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_26_6_0 INVX1_3/gnd DFFSR_23/S FILL
XFILL_12_DFFSR_221 AND2X2_38/B DFFSR_59/S FILL
XFILL_22_DFFPOSX1_44 OR2X2_2/gnd DFFSR_216/S FILL
XDFFSR_111 DFFSR_119/D CLKBUF1_5/Y DFFSR_35/R DFFSR_8/S AOI22X1_7/B DFFSR_8/gnd DFFSR_8/S
+ DFFSR
XFILL_4_DFFSR_108 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_6_NAND3X1_247 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_1_BUFX2_38 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_1_OAI22X1_1 INVX1_1/gnd DFFSR_53/S FILL
XFILL_45_DFFSR_139 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_8_DFFSR_215 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_35_DFFSR_142 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_49_DFFSR_246 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_11_DFFSR_4 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_25_DFFSR_145 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_39_DFFSR_249 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_1_INVX1_192 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_38_DFFSR_60 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_49_DFFSR_20 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_15_DFFSR_148 INVX1_67/gnd DFFSR_175/S FILL
XFILL_7_NAND3X1_181 INVX1_39/gnd DFFSR_54/S FILL
XFILL_29_DFFSR_252 AND2X2_38/B DFFSR_23/S FILL
XFILL_0_NAND2X1_162 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_19_DFFSR_255 OR2X2_4/gnd DFFSR_32/S FILL
XDFFSR_57 INVX1_2/A DFFSR_57/CLK DFFSR_3/R DFFSR_6/S DFFSR_57/D BUFX2_79/A DFFSR_6/S
+ DFFSR
XFILL_5_DFFSR_17 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_22_DFFSR_10 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_11_DFFSR_50 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_0_NOR2X1_27 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_8_NAND3X1_115 BUFX2_79/A DFFSR_7/S FILL
XINVX1_122 NOR3X1_1/A DFFSR_1/gnd INVX1_122/Y DFFSR_1/S INVX1
XFILL_1_DFFSR_145 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_12_DFFPOSX1_19 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_42_DFFSR_176 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_4_INVX1_119 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_46_DFFSR_67 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_5_DFFSR_252 AND2X2_38/B DFFSR_23/S FILL
XFILL_32_DFFSR_179 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_36_1_0 BUFX2_99/A DFFSR_92/S FILL
XFILL_22_DFFSR_182 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_30_DFFSR_17 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_2_DFFSR_64 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_2_INVX1_11 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_19_DFFSR_57 BUFX2_79/A DFFSR_6/S FILL
XFILL_12_DFFSR_185 INVX1_39/gnd DFFSR_54/S FILL
XFILL_6_BUFX2_92 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_34_3_1 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_9_OAI21X1_9 INVX1_67/gnd DFFSR_201/S FILL
XFILL_20_CLKBUF1_47 BUFX2_98/A DFFSR_32/S FILL
XFILL_6_NAND3X1_211 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_45_DFFSR_103 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_32_5_2 INVX1_1/gnd DFFSR_97/S FILL
XFILL_2_DFFPOSX1_30 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_8_DFFSR_179 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_35_DFFSR_106 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_49_DFFSR_210 BUFX2_98/A DFFSR_6/S FILL
XAND2X2_26 AND2X2_26/A AND2X2_26/B INVX1_1/gnd AND2X2_26/Y DFFSR_97/S AND2X2
XFILL_25_DFFSR_109 DFFSR_4/gnd DFFSR_4/S FILL
XNAND3X1_247 BUFX2_8/Y OR2X2_1/A NOR3X1_1/A NOR3X1_6/gnd NOR3X1_6/C DFFSR_79/S NAND3X1
XFILL_38_DFFSR_24 BUFX2_98/A DFFSR_6/S FILL
XFILL_39_DFFSR_213 INVX1_3/gnd DFFSR_23/S FILL
XFILL_1_INVX1_156 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_27_DFFSR_64 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_4_AND2X2_23 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_15_DFFSR_112 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_7_NAND3X1_145 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_29_DFFSR_216 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_11_DFFPOSX1_49 BUFX2_99/A DFFSR_92/S FILL
XFILL_19_DFFSR_219 INVX1_67/gnd DFFSR_175/S FILL
XFILL_0_NAND2X1_126 OR2X2_2/gnd DFFSR_175/S FILL
XDFFSR_21 INVX1_35/A DFFSR_82/CLK DFFSR_5/R DFFSR_5/S INVX1_36/A DFFSR_5/gnd DFFSR_5/S
+ DFFSR
XFILL_11_DFFSR_14 INVX1_1/gnd DFFSR_53/S FILL
XFILL_1_DFFSR_109 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_21_DFFPOSX1_38 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_42_DFFSR_140 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_46_DFFSR_31 BUFX2_79/A DFFSR_6/S FILL
XFILL_35_DFFSR_71 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_5_DFFSR_216 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_32_DFFSR_143 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_5_NAND3X1_241 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_46_DFFSR_247 BUFX2_99/A DFFSR_7/S FILL
XFILL_22_DFFSR_146 BUFX2_79/A DFFSR_7/S FILL
XFILL_2_DFFSR_28 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_36_DFFSR_250 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_19_DFFSR_21 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_12_DFFSR_149 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_6_BUFX2_56 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_26_DFFSR_253 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_42_0_2 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_16_DFFSR_256 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_1_NOR2X1_9 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_6_NAND3X1_175 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_20_CLKBUF1_11 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_19_CLKBUF1_14 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_8_DFFSR_143 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_43_DFFSR_78 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_49_DFFSR_174 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_18_CLKBUF1_17 BUFX2_8/gnd DFFSR_81/S FILL
XNAND3X1_211 OAI21X1_71/Y INVX1_164/Y OAI21X1_72/Y DFFSR_1/gnd NAND3X1_215/B DFFSR_81/S
+ NAND3X1
XFILL_17_CLKBUF1_20 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_39_DFFSR_177 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_1_INVX1_120 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_27_DFFSR_28 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_16_DFFSR_68 BUFX2_98/A DFFSR_6/S FILL
XFILL_7_NAND3X1_109 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_2_DFFSR_253 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_16_CLKBUF1_23 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_29_DFFSR_180 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_11_DFFPOSX1_13 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_19_DFFSR_183 INVX1_67/gnd DFFSR_175/S FILL
XFILL_15_CLKBUF1_26 INVX1_1/gnd DFFSR_53/S FILL
XNOR2X1_65 NOR2X1_66/B NOR2X1_65/B DFFSR_34/gnd NOR2X1_65/Y DFFSR_1/S NOR2X1
XFILL_14_CLKBUF1_29 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_3_XOR2X1_5 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_4_NOR2X1_62 INVX1_67/gnd DFFSR_201/S FILL
XFILL_23_DFFSR_7 BUFX2_79/A DFFSR_7/S FILL
XFILL_13_CLKBUF1_32 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_12_CLKBUF1_35 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_42_DFFSR_104 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_35_DFFSR_35 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_11_CLKBUF1_38 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_7_DFFSR_82 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_24_DFFSR_75 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_5_DFFSR_180 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_32_DFFSR_107 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_46_DFFSR_211 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_10_CLKBUF1_41 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_5_NAND3X1_205 INVX1_1/gnd DFFSR_53/S FILL
XFILL_22_DFFSR_110 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_36_DFFSR_214 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_1_DFFPOSX1_24 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_1_AND2X2_24 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_6_BUFX2_20 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_12_DFFSR_113 BUFX2_99/A DFFSR_92/S FILL
XFILL_5_NAND2X1_1 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_26_DFFSR_217 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_9_CLKBUF1_44 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_16_DFFSR_220 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_8_CLKBUF1_47 BUFX2_98/A DFFSR_32/S FILL
XFILL_44_DFFSR_3 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_6_NAND3X1_139 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_10_DFFPOSX1_43 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_4_INVX1_76 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_32_DFFSR_82 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_43_DFFSR_42 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_8_DFFSR_107 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_49_DFFSR_138 BUFX2_8/gnd DFFSR_81/S FILL
XNAND3X1_175 INVX1_135/A AND2X2_33/B NOR2X1_70/B NOR3X1_6/gnd NAND3X1_176/C DFFSR_91/S
+ NAND3X1
XFILL_39_DFFSR_141 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_16_DFFSR_32 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_22_3 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_2_DFFSR_217 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_3_BUFX2_67 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_29_DFFSR_144 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_33_6_0 INVX1_1/gnd DFFSR_53/S FILL
XFILL_43_DFFSR_248 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_20_DFFPOSX1_32 INVX1_67/gnd DFFSR_201/S FILL
XFILL_19_DFFSR_147 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_33_DFFSR_251 BUFX2_7/gnd DFFSR_151/S FILL
XNOR2X1_29 NOR2X1_29/A NOR2X1_29/B DFFSR_28/gnd NOR2X1_29/Y DFFSR_3/S NOR2X1
XFILL_23_DFFSR_254 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_4_NAND3X1_235 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_40_DFFSR_89 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_4_NOR2X1_26 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_13_DFFSR_257 INVX1_39/gnd DFFSR_34/S FILL
XFILL_24_DFFSR_39 INVX1_3/gnd DFFSR_79/S FILL
XFILL_7_DFFSR_46 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_13_DFFSR_79 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_5_DFFSR_144 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_46_DFFSR_175 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_5_NAND3X1_169 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_9_DFFSR_251 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_36_DFFSR_178 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_26_DFFSR_181 INVX1_3/gnd DFFSR_79/S FILL
XFILL_48_DFFSR_96 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_16_DFFSR_184 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_10_DFFSR_1 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_8_CLKBUF1_11 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_6_NAND3X1_103 AND2X2_38/B DFFSR_23/S FILL
XFILL_7_CLKBUF1_14 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_4_INVX1_40 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_4_DFFSR_93 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_21_DFFSR_86 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_32_DFFSR_46 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_1_NOR2X1_63 INVX1_3/gnd DFFSR_23/S FILL
XFILL_6_CLKBUF1_17 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_49_DFFSR_102 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_43_1_0 OR2X2_4/gnd DFFSR_3/S FILL
XNAND3X1_139 AND2X2_35/A INVX1_135/A AND2X2_29/Y BUFX2_8/gnd OAI21X1_30/C DFFSR_51/S
+ NAND3X1
XFILL_5_CLKBUF1_20 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_39_DFFSR_105 INVX1_1/gnd DFFSR_53/S FILL
XCLKBUF1_17 BUFX2_4/Y BUFX2_8/gnd CLKBUF1_17/Y DFFSR_81/S CLKBUF1
XFILL_5_7 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_4_CLKBUF1_23 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_2_DFFSR_181 INVX1_3/gnd DFFSR_79/S FILL
XFILL_3_BUFX2_31 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_29_DFFSR_108 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_43_DFFSR_212 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_3_CLKBUF1_26 INVX1_1/gnd DFFSR_53/S FILL
XFILL_8_AND2X2_22 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_19_DFFSR_111 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_41_3_1 BUFX2_98/A DFFSR_32/S FILL
XFILL_2_CLKBUF1_29 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_33_DFFSR_215 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_2_NAND2X1_2 BUFX2_99/A DFFSR_7/S FILL
XFILL_23_DFFSR_218 BUFX2_98/A DFFSR_32/S FILL
XFILL_4_NAND3X1_199 INVX1_1/gnd DFFSR_97/S FILL
XFILL_1_CLKBUF1_32 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_1_INVX1_87 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_40_DFFSR_53 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_29_DFFSR_93 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_39_5_2 BUFX2_79/A DFFSR_6/S FILL
XFILL_0_CLKBUF1_35 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_13_DFFSR_221 AND2X2_38/B DFFSR_59/S FILL
XFILL_0_DFFPOSX1_18 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_7_DFFSR_10 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_13_DFFSR_43 BUFX2_98/A DFFSR_6/S FILL
XFILL_5_DFFSR_108 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_0_BUFX2_78 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_2_OAI22X1_1 INVX1_1/gnd DFFSR_53/S FILL
XFILL_9_OR2X2_6 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_46_DFFSR_139 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_5_NAND3X1_133 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_9_DFFSR_215 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_36_DFFSR_142 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_50_DFFSR_246 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_26_DFFSR_145 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_40_DFFSR_249 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_2_INVX1_192 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_48_DFFSR_60 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_16_DFFSR_148 INVX1_67/gnd DFFSR_175/S FILL
XFILL_44_3 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_30_DFFSR_252 AND2X2_38/B DFFSR_23/S FILL
XFILL_20_DFFSR_255 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_4_DFFSR_57 BUFX2_79/A DFFSR_6/S FILL
XFILL_32_DFFSR_10 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_21_DFFSR_50 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_10_DFFSR_90 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_19_DFFPOSX1_26 AND2X2_38/B DFFSR_23/S FILL
XFILL_1_NOR2X1_27 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_10_DFFSR_258 DFFSR_5/gnd DFFSR_5/S FILL
XNAND3X1_103 NAND3X1_103/A NAND3X1_103/B AOI22X1_13/Y AND2X2_38/B NOR2X1_49/B DFFSR_23/S
+ NAND3X1
XFILL_3_NAND3X1_229 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_2_DFFSR_145 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_43_DFFSR_176 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_6_DFFSR_252 AND2X2_38/B DFFSR_23/S FILL
XFILL_49_0_2 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_33_DFFSR_179 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_23_DFFSR_182 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_4_NAND3X1_163 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_40_DFFSR_17 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_1_INVX1_51 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_29_DFFSR_57 BUFX2_79/A DFFSR_6/S FILL
XFILL_18_DFFSR_97 INVX1_1/gnd DFFSR_97/S FILL
XFILL_13_DFFSR_185 INVX1_39/gnd DFFSR_54/S FILL
XFILL_9_DFFPOSX1_37 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_0_BUFX2_42 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_46_DFFSR_103 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_9_DFFSR_179 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_36_DFFSR_106 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_50_DFFSR_210 BUFX2_98/A DFFSR_6/S FILL
XFILL_26_DFFSR_109 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_40_DFFSR_213 INVX1_3/gnd DFFSR_23/S FILL
XFILL_2_INVX1_156 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_37_DFFSR_64 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_48_DFFSR_24 BUFX2_98/A DFFSR_6/S FILL
XFILL_5_AND2X2_23 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_16_DFFSR_112 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_30_DFFSR_216 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_15_1_1 INVX1_39/gnd DFFSR_34/S FILL
XFILL_20_DFFSR_219 INVX1_67/gnd DFFSR_175/S FILL
XFILL_4_DFFSR_21 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_21_DFFSR_14 INVX1_1/gnd DFFSR_53/S FILL
XFILL_10_DFFSR_54 INVX1_39/gnd DFFSR_54/S FILL
XFILL_5_OAI21X1_115 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_10_DFFSR_222 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_13_3_2 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_3_NAND3X1_193 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_2_DFFSR_109 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_3_NOR2X1_2 INVX1_1/gnd DFFSR_97/S FILL
XFILL_22_DFFSR_4 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_43_DFFSR_140 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_45_DFFSR_71 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_6_DFFSR_216 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_33_DFFSR_143 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_47_DFFSR_247 BUFX2_99/A DFFSR_7/S FILL
XFILL_23_DFFSR_146 BUFX2_79/A DFFSR_7/S FILL
XFILL_4_NAND3X1_127 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_37_DFFSR_250 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_29_DFFSR_21 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_1_INVX1_15 BUFX2_98/A DFFSR_32/S FILL
XFILL_1_DFFSR_68 BUFX2_98/A DFFSR_6/S FILL
XFILL_18_DFFSR_61 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_13_DFFSR_149 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_5_BUFX2_96 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_6_BUFX2_5 AND2X2_38/B DFFSR_59/S FILL
XFILL_27_DFFSR_253 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_6_NAND2X1_163 INVX1_67/gnd DFFSR_201/S FILL
XFILL_17_DFFSR_256 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_49_8 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_9_DFFSR_143 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_40_6_0 BUFX2_98/A DFFSR_6/S FILL
XFILL_18_DFFPOSX1_20 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_50_DFFSR_174 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_19_DFFPOSX1_2 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_40_DFFSR_177 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_2_INVX1_120 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_37_DFFSR_28 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_26_DFFSR_68 BUFX2_98/A DFFSR_6/S FILL
XFILL_9_DFFSR_75 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_2_NAND3X1_223 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_18_DFFPOSX1_5 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_3_DFFSR_253 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_30_DFFSR_180 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_17_DFFPOSX1_8 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_20_DFFSR_183 INVX1_67/gnd DFFSR_175/S FILL
XFILL_10_DFFSR_18 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_10_DFFSR_186 BUFX2_99/A DFFSR_92/S FILL
XFILL_5_NOR2X1_62 INVX1_67/gnd DFFSR_201/S FILL
XFILL_3_NAND3X1_157 INVX1_3/gnd DFFSR_23/S FILL
XFILL_43_DFFSR_104 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_8_DFFPOSX1_31 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_45_DFFSR_35 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_34_DFFSR_75 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_6_DFFSR_180 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_33_DFFSR_107 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_47_DFFSR_211 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_23_DFFSR_110 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_37_DFFSR_214 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_1_DFFSR_32 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_18_DFFSR_25 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_2_AND2X2_24 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_13_DFFSR_113 BUFX2_99/A DFFSR_92/S FILL
XFILL_5_BUFX2_60 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_6_NAND2X1_1 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_27_DFFSR_217 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_17_DFFPOSX1_50 INVX1_1/gnd DFFSR_53/S FILL
XFILL_10_OAI22X1_6 BUFX2_98/A DFFSR_32/S FILL
XFILL_6_NAND2X1_127 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_17_DFFSR_220 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_50_1_0 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_9_NOR3X1_6 NOR3X1_6/gnd DFFSR_79/S FILL
XXOR2X1_2 XOR2X1_2/A XOR2X1_2/B OR2X2_2/gnd OR2X2_2/A DFFSR_175/S XOR2X1
XFILL_42_DFFSR_82 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_9_DFFSR_107 OR2X2_6/gnd DFFSR_92/S FILL
XNAND2X1_163 DFFSR_175/S NAND2X1_163/B INVX1_67/gnd AOI21X1_57/B DFFSR_201/S NAND2X1
XFILL_48_3_1 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_50_DFFSR_138 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_4_OAI21X1_109 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_27_DFFPOSX1_39 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_8_AOI21X1_55 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_40_DFFSR_141 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_7_AOI21X1_58 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_15_DFFSR_72 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_26_DFFSR_32 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_9_DFFSR_39 INVX1_3/gnd DFFSR_79/S FILL
XFILL_2_NAND3X1_187 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_3_DFFSR_217 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_46_5_2 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_30_DFFSR_144 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_6_AOI21X1_61 AND2X2_38/B DFFSR_59/S FILL
XFILL_44_DFFSR_248 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_20_DFFSR_147 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_5_AOI21X1_64 AND2X2_38/B DFFSR_59/S FILL
XFILL_34_DFFSR_251 BUFX2_7/gnd DFFSR_151/S FILL
XAOI21X1_61 OR2X2_1/B OR2X2_1/A AOI21X1_61/C AND2X2_38/B AOI21X1_61/Y DFFSR_59/S AOI21X1
XFILL_10_DFFSR_150 AND2X2_38/B DFFSR_23/S FILL
XFILL_4_AOI21X1_67 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_2_XOR2X1_9 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_24_DFFSR_254 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_50_DFFSR_89 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_5_NOR2X1_26 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_3_NAND3X1_121 INVX1_1/gnd DFFSR_97/S FILL
XFILL_3_AOI21X1_70 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_14_DFFSR_257 INVX1_39/gnd DFFSR_34/S FILL
XFILL_6_DFFSR_86 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_5_NAND2X1_157 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_23_DFFSR_79 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_34_DFFSR_39 INVX1_3/gnd DFFSR_79/S FILL
XFILL_6_DFFSR_144 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_14_4_0 INVX1_39/gnd DFFSR_54/S FILL
XFILL_47_DFFSR_175 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_37_DFFSR_178 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_8_OR2X2_3 OR2X2_3/gnd DFFSR_4/S FILL
XBUFX2_64 BUFX2_60/A DFFSR_62/gnd BUFX2_64/Y DFFSR_62/S BUFX2
XFILL_5_BUFX2_24 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_0_DFFSR_254 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_27_DFFSR_181 INVX1_3/gnd DFFSR_79/S FILL
XFILL_12_6_1 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_17_DFFPOSX1_14 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_17_DFFSR_184 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_34_DFFSR_7 BUFX2_79/A DFFSR_7/S FILL
XFILL_15_NOR3X1_3 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_1_NAND3X1_217 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_31_DFFSR_86 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_3_INVX1_80 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_42_DFFSR_46 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_2_NOR2X1_63 INVX1_3/gnd DFFSR_23/S FILL
XNAND2X1_127 BUFX2_55/Y INVX1_148/A OR2X2_1/gnd OAI21X1_96/C DFFSR_51/S NAND2X1
XFILL_50_DFFSR_102 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_7_DFFPOSX1_2 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_8_AOI21X1_19 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_40_DFFSR_105 INVX1_1/gnd DFFSR_53/S FILL
XFILL_6_DFFPOSX1_5 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_9_4 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_15_DFFSR_36 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_7_AOI21X1_22 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_2_NAND3X1_151 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_3_DFFSR_181 INVX1_3/gnd DFFSR_79/S FILL
XFILL_2_BUFX2_71 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_30_DFFSR_108 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_5_DFFPOSX1_8 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_6_AOI21X1_25 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_44_DFFSR_212 OR2X2_2/gnd DFFSR_175/S FILL
XDFFPOSX1_5 DFFPOSX1_5/Q CLKBUF1_44/Y NOR2X1_60/Y OR2X2_2/gnd DFFSR_216/S DFFPOSX1
XFILL_20_DFFSR_111 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_7_DFFPOSX1_25 BUFX2_79/A DFFSR_6/S FILL
XFILL_5_AOI21X1_28 AND2X2_38/B DFFSR_23/S FILL
XFILL_34_DFFSR_215 DFFSR_34/gnd DFFSR_1/S FILL
XAOI21X1_25 AOI21X1_25/A AOI21X1_25/B NAND2X1_79/B DFFSR_62/gnd AOI21X1_25/Y DFFSR_208/S
+ AOI21X1
XFILL_3_NAND2X1_2 BUFX2_99/A DFFSR_7/S FILL
XFILL_10_DFFSR_114 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_24_DFFSR_218 BUFX2_98/A DFFSR_32/S FILL
XFILL_4_AOI21X1_31 INVX1_39/gnd DFFSR_34/S FILL
XFILL_50_DFFSR_53 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_39_DFFSR_93 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_3_AOI21X1_34 INVX1_39/gnd DFFSR_34/S FILL
XFILL_14_DFFSR_221 AND2X2_38/B DFFSR_59/S FILL
XFILL_16_DFFPOSX1_44 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_2_AOI21X1_37 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_0_AND2X2_2 BUFX2_99/A DFFSR_7/S FILL
XFILL_6_DFFSR_50 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_5_NAND2X1_121 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_23_DFFSR_43 BUFX2_98/A DFFSR_6/S FILL
XFILL_6_DFFSR_108 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_12_DFFSR_83 INVX1_3/gnd DFFSR_79/S FILL
XFILL_1_AOI21X1_40 INVX1_39/gnd DFFSR_54/S FILL
XFILL_3_OAI22X1_1 INVX1_1/gnd DFFSR_53/S FILL
XFILL_0_NAND3X1_247 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_47_DFFSR_139 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_0_AOI21X1_43 INVX1_3/gnd DFFSR_79/S FILL
XFILL_22_1_1 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_37_DFFSR_142 XOR2X1_1/gnd DFFSR_151/S FILL
XBUFX2_28 BUFX2_27/A DFFSR_46/gnd BUFX2_28/Y DFFSR_62/S BUFX2
XFILL_4_0_0 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_0_DFFSR_218 BUFX2_98/A DFFSR_32/S FILL
XFILL_27_DFFSR_145 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_3_OAI21X1_103 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_41_DFFSR_249 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_3_INVX1_192 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_26_DFFPOSX1_33 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_31_5 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_20_3_2 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_17_DFFSR_148 INVX1_67/gnd DFFSR_175/S FILL
XFILL_8_OAI21X1_67 INVX1_1/gnd DFFSR_97/S FILL
XFILL_31_DFFSR_252 AND2X2_38/B DFFSR_23/S FILL
XFILL_1_NAND3X1_181 INVX1_39/gnd DFFSR_54/S FILL
XFILL_2_2_1 INVX1_67/gnd DFFSR_201/S FILL
XFILL_8_AND2X2_9 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_7_OAI21X1_70 INVX1_3/gnd DFFSR_23/S FILL
XFILL_6_NAND2X1_88 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_21_DFFSR_255 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_42_DFFSR_10 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_31_DFFSR_50 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_3_INVX1_44 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_3_DFFSR_97 INVX1_1/gnd DFFSR_97/S FILL
XFILL_2_NOR2X1_27 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_20_DFFSR_90 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_5_NAND2X1_91 INVX1_39/gnd DFFSR_54/S FILL
XFILL_6_OAI21X1_73 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_11_DFFSR_258 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_0_4_2 BUFX2_72/gnd DFFSR_276/S FILL
XNAND2X1_88 AOI22X1_23/A AOI22X1_23/B DFFSR_34/gnd OAI21X1_58/C DFFSR_1/S NAND2X1
XFILL_4_NAND2X1_94 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_5_OAI21X1_76 INVX1_1/gnd DFFSR_53/S FILL
XOAI21X1_73 OAI21X1_73/A OAI21X1_73/B AOI21X1_22/C DFFSR_46/gnd AOI21X1_32/A DFFSR_54/S
+ OAI21X1
XFILL_3_DFFSR_145 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_2_NAND3X1_115 BUFX2_79/A DFFSR_7/S FILL
XFILL_4_OAI21X1_79 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_3_NAND2X1_97 INVX1_1/gnd DFFSR_97/S FILL
XFILL_2_BUFX2_35 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_44_DFFSR_176 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_3_OAI21X1_82 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_7_DFFSR_252 AND2X2_38/B DFFSR_23/S FILL
XFILL_34_DFFSR_179 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_4_NAND2X1_151 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_2_OAI21X1_85 INVX1_39/gnd DFFSR_54/S FILL
XFILL_21_DFFSR_1 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_24_DFFSR_182 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_50_DFFSR_17 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_1_OAI21X1_88 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_39_DFFSR_57 BUFX2_79/A DFFSR_6/S FILL
XFILL_28_DFFSR_97 INVX1_1/gnd DFFSR_97/S FILL
XFILL_0_INVX1_91 AND2X2_38/B DFFSR_23/S FILL
XFILL_47_6_0 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_14_DFFSR_185 INVX1_39/gnd DFFSR_54/S FILL
XFILL_0_OAI21X1_91 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_6_DFFSR_14 INVX1_1/gnd DFFSR_53/S FILL
XFILL_12_DFFSR_47 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_5_BUFX2_2 OR2X2_4/gnd DFFSR_32/S FILL
XBUFX2_6 BUFX2_3/A BUFX2_79/A BUFX2_6/Y DFFSR_6/S BUFX2
XFILL_0_NAND3X1_211 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_47_DFFSR_103 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_37_DFFSR_106 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_0_DFFSR_182 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_27_DFFSR_109 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_9_OAI21X1_28 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_41_DFFSR_213 INVX1_3/gnd DFFSR_23/S FILL
XFILL_3_INVX1_156 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_47_DFFSR_64 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_6_AND2X2_23 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_17_DFFSR_112 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_31_DFFSR_216 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_8_OAI21X1_31 AND2X2_38/B DFFSR_23/S FILL
XFILL_1_NAND3X1_145 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_0_NAND2X1_3 BUFX2_99/A DFFSR_7/S FILL
XFILL_7_OAI21X1_34 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_6_NAND2X1_52 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_21_DFFSR_219 INVX1_67/gnd DFFSR_175/S FILL
XFILL_3_DFFSR_61 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_31_DFFSR_14 INVX1_1/gnd DFFSR_53/S FILL
XFILL_20_DFFSR_54 INVX1_39/gnd DFFSR_54/S FILL
XFILL_6_DFFPOSX1_19 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_6_OAI21X1_37 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_5_NAND2X1_55 INVX1_39/gnd DFFSR_34/S FILL
XFILL_11_DFFSR_222 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_3_NAND2X1_181 BUFX2_99/A DFFSR_92/S FILL
XNAND2X1_52 DFFSR_176/D AND2X2_18/Y OR2X2_6/gnd NAND2X1_52/Y DFFSR_53/S NAND2X1
XFILL_4_NAND2X1_58 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_5_OAI21X1_40 DFFSR_34/gnd DFFSR_1/S FILL
XOAI21X1_37 INVX1_143/A NAND2X1_71/Y OAI21X1_37/C DFFSR_1/gnd INVX1_152/A DFFSR_81/S
+ OAI21X1
XFILL_3_DFFSR_109 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_3_NAND2X1_61 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_4_OAI21X1_43 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_0_OAI22X1_2 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_44_DFFSR_140 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_15_DFFPOSX1_38 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_3_OAI21X1_46 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_2_NAND2X1_64 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_7_DFFSR_216 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_34_DFFSR_143 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_4_NAND2X1_115 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_1_NAND2X1_67 AND2X2_38/B DFFSR_59/S FILL
XFILL_2_OAI21X1_49 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_48_DFFSR_247 BUFX2_99/A DFFSR_7/S FILL
XFILL_11_AOI22X1_15 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_24_DFFSR_146 BUFX2_79/A DFFSR_7/S FILL
XFILL_0_NAND2X1_70 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_38_DFFSR_250 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_1_OAI21X1_52 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_28_DFFSR_61 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_0_INVX1_55 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_39_DFFSR_21 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_10_AOI22X1_18 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_0_INVX1_193 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_14_DFFSR_149 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_28_DFFSR_253 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_0_OAI21X1_55 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_53_5 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_18_DFFSR_256 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_25_DFFPOSX1_27 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_9_AOI22X1_21 AND2X2_38/B DFFSR_59/S FILL
XFILL_12_DFFSR_11 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_0_NAND3X1_175 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_8_AOI22X1_24 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_53_5_2 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_7_AOI22X1_27 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_5_DFFPOSX1_49 BUFX2_99/A DFFSR_92/S FILL
XDFFSR_256 BUFX2_97/A DFFSR_85/CLK BUFX2_65/Y DFFSR_60/S INVX1_117/A DFFSR_8/gnd DFFSR_60/S
+ DFFSR
XFILL_0_DFFSR_146 BUFX2_79/A DFFSR_7/S FILL
XFILL_41_DFFSR_177 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_3_INVX1_120 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_47_DFFSR_28 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_36_DFFSR_68 BUFX2_98/A DFFSR_6/S FILL
XFILL_4_DFFSR_253 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_31_DFFSR_180 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_1_NAND3X1_109 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_6_NAND2X1_16 BUFX2_79/A DFFSR_7/S FILL
XFILL_21_DFFSR_183 INVX1_67/gnd DFFSR_175/S FILL
XFILL_3_DFFSR_25 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_20_DFFSR_18 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_3_NAND2X1_145 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_5_NAND2X1_19 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_11_DFFSR_186 BUFX2_99/A DFFSR_92/S FILL
XNAND2X1_16 DFFSR_43/D AND2X2_5/Y BUFX2_79/A NAND3X1_20/A DFFSR_7/S NAND2X1
XFILL_4_NAND2X1_22 BUFX2_99/A DFFSR_7/S FILL
XFILL_21_4_0 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_6_NOR2X1_62 INVX1_67/gnd DFFSR_201/S FILL
XFILL_2_NOR2X1_6 BUFX2_98/A DFFSR_6/S FILL
XFILL_3_NAND2X1_25 BUFX2_99/A DFFSR_7/S FILL
XDFFPOSX1_19 INVX1_162/A CLKBUF1_44/Y OAI21X1_57/Y DFFSR_34/gnd DFFSR_1/S DFFPOSX1
XFILL_44_DFFSR_104 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_12_DFFSR_8 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_3_OAI21X1_10 BUFX2_79/A DFFSR_7/S FILL
XFILL_2_NAND2X1_28 AND2X2_38/B DFFSR_59/S FILL
XFILL_19_6_1 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_44_DFFSR_75 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_7_DFFSR_180 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_34_DFFSR_107 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_9_NAND3X1_84 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_1_NAND2X1_31 INVX1_3/gnd DFFSR_23/S FILL
XFILL_2_OAI21X1_13 INVX1_39/gnd DFFSR_54/S FILL
XFILL_1_5_0 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_48_DFFSR_211 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_24_DFFSR_110 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_0_NAND2X1_34 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_8_NAND3X1_87 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_38_DFFSR_214 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_1_OAI21X1_16 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_0_INVX1_19 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_0_INVX1_157 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_0_DFFSR_72 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_28_DFFSR_25 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_17_DFFSR_65 BUFX2_79/A DFFSR_7/S FILL
XFILL_3_AND2X2_24 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_14_DFFSR_113 BUFX2_99/A DFFSR_92/S FILL
XFILL_7_NAND3X1_90 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_28_DFFSR_217 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_0_OAI21X1_19 BUFX2_98/A DFFSR_32/S FILL
XFILL_11_OAI22X1_6 BUFX2_98/A DFFSR_32/S FILL
XFILL_6_NAND3X1_93 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_18_DFFSR_220 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_5_NAND3X1_96 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_0_NAND3X1_139 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_4_XOR2X1_2 OR2X2_2/gnd DFFSR_175/S FILL
XNAND3X1_93 DFFSR_196/D BUFX2_34/Y BUFX2_23/Y XOR2X1_1/gnd NAND3X1_93/Y DFFSR_208/S
+ NAND3X1
XFILL_4_NAND3X1_99 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_9_NAND3X1_194 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_33_DFFSR_4 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_5_DFFPOSX1_13 BUFX2_8/gnd DFFSR_81/S FILL
XDFFSR_220 DFFSR_220/Q CLKBUF1_31/Y BUFX2_60/Y DFFSR_151/S INVX1_85/A BUFX2_7/gnd
+ DFFSR_151/S DFFSR
XFILL_0_DFFSR_110 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_2_NAND2X1_175 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_13_2 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_41_DFFSR_141 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_36_DFFSR_32 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_8_DFFSR_79 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_25_DFFSR_72 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_4_DFFSR_217 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_31_DFFSR_144 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_45_DFFSR_248 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_21_DFFSR_147 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_14_DFFPOSX1_32 INVX1_67/gnd DFFSR_201/S FILL
XFILL_35_DFFSR_251 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_3_NAND2X1_109 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_11_DFFSR_150 AND2X2_38/B DFFSR_23/S FILL
XFILL_25_DFFSR_254 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_6_NOR2X1_26 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_29_1_1 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_15_DFFSR_257 INVX1_39/gnd DFFSR_34/S FILL
XFILL_0_NOR3X1_3 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_10_OAI22X1_30 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_0_AOI22X1_12 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_33_DFFSR_79 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_44_DFFSR_39 INVX1_3/gnd DFFSR_79/S FILL
XFILL_7_DFFSR_144 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_24_DFFPOSX1_21 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_9_NAND3X1_48 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_27_3_2 INVX1_3/gnd DFFSR_79/S FILL
XFILL_48_DFFSR_175 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_8_NAND3X1_51 BUFX2_99/A DFFSR_7/S FILL
XFILL_9_OAI22X1_33 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_9_2_1 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_38_DFFSR_178 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_0_INVX1_121 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_8_NAND3X1_224 INVX1_39/gnd DFFSR_54/S FILL
XFILL_17_DFFSR_29 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_0_DFFSR_36 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_8_OAI22X1_36 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_7_NAND3X1_54 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_1_DFFSR_254 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_4_BUFX2_64 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_28_DFFSR_181 INVX1_3/gnd DFFSR_79/S FILL
XFILL_4_DFFPOSX1_43 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_6_NAND3X1_57 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_7_OAI22X1_39 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_7_4_2 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_18_DFFSR_184 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_5_NAND3X1_60 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_6_OAI22X1_42 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_0_NAND3X1_103 AND2X2_38/B DFFSR_23/S FILL
XNAND3X1_57 DFFSR_48/Q BUFX2_17/Y BUFX2_12/Y DFFSR_8/gnd NAND3X1_60/B DFFSR_60/S NAND3X1
XFILL_5_OAI22X1_45 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_4_NAND3X1_63 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_41_DFFSR_86 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_3_NOR2X1_63 INVX1_3/gnd DFFSR_23/S FILL
XOAI22X1_42 INVX1_101/Y OAI22X1_45/B INVX1_102/Y OAI22X1_45/D BUFX2_8/gnd NOR2X1_51/A
+ DFFSR_51/S OAI22X1
XFILL_3_NAND3X1_66 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_4_OAI22X1_48 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_2_NAND2X1_139 INVX1_1/gnd DFFSR_97/S FILL
XDFFSR_184 DFFSR_144/D CLKBUF1_22/Y BUFX2_70/Y DFFSR_51/S DFFSR_184/D OR2X2_1/gnd
+ DFFSR_51/S DFFSR
XFILL_2_NAND3X1_69 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_41_DFFSR_105 INVX1_1/gnd DFFSR_53/S FILL
XFILL_3_OAI22X1_51 INVX1_39/gnd DFFSR_54/S FILL
XFILL_8_DFFSR_43 BUFX2_98/A DFFSR_6/S FILL
XFILL_25_DFFSR_36 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_14_DFFSR_76 BUFX2_79/A DFFSR_7/S FILL
XFILL_4_DFFSR_181 INVX1_3/gnd DFFSR_79/S FILL
XFILL_31_DFFSR_108 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_1_NAND3X1_72 INVX1_39/gnd DFFSR_34/S FILL
XFILL_45_DFFSR_212 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_54_6_0 DFFSR_5/gnd DFFSR_5/S FILL
XNAND2X1_5 NOR2X1_4/Y AND2X2_2/Y OR2X2_4/gnd OAI22X1_6/D DFFSR_3/S NAND2X1
XFILL_21_DFFSR_111 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_0_NAND3X1_75 BUFX2_79/A DFFSR_7/S FILL
XFILL_35_DFFSR_215 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_0_AND2X2_25 INVX1_39/gnd DFFSR_54/S FILL
XFILL_4_NAND2X1_2 BUFX2_99/A DFFSR_7/S FILL
XFILL_11_DFFSR_114 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_25_DFFSR_218 BUFX2_98/A DFFSR_32/S FILL
XFILL_0_DFFSR_7 BUFX2_79/A DFFSR_7/S FILL
XFILL_49_DFFSR_93 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_15_DFFSR_221 AND2X2_38/B DFFSR_59/S FILL
XOAI22X1_4 INVX1_10/Y OAI22X1_7/B INVX1_11/Y OAI22X1_7/D OR2X2_3/gnd NOR2X1_9/B DFFSR_4/S
+ OAI22X1
XINVX1_77 INVX1_77/A DFFSR_1/gnd INVX1_77/Y DFFSR_81/S INVX1
XFILL_5_DFFSR_90 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_33_DFFSR_43 BUFX2_98/A DFFSR_6/S FILL
XFILL_7_DFFSR_108 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_22_DFFSR_83 INVX1_3/gnd DFFSR_79/S FILL
XFILL_4_OAI22X1_1 INVX1_1/gnd DFFSR_53/S FILL
XFILL_48_DFFSR_139 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_8_NAND3X1_15 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_8_NAND3X1_188 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_38_DFFSR_142 XOR2X1_1/gnd DFFSR_151/S FILL
XINVX1_195 INVX1_195/A DFFSR_46/gnd INVX1_195/Y DFFSR_54/S INVX1
XFILL_1_DFFSR_218 BUFX2_98/A DFFSR_32/S FILL
XFILL_7_NAND3X1_18 BUFX2_79/A DFFSR_7/S FILL
XFILL_4_BUFX2_28 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_28_DFFSR_145 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_42_DFFSR_249 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_1_NAND2X1_169 INVX1_1/gnd DFFSR_53/S FILL
XFILL_6_NAND3X1_21 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_18_DFFSR_148 INVX1_67/gnd DFFSR_175/S FILL
XFILL_32_DFFSR_252 AND2X2_38/B DFFSR_23/S FILL
XFILL_5_NAND3X1_24 INVX1_1/gnd DFFSR_97/S FILL
XNAND3X1_21 DFFSR_67/D BUFX2_22/Y BUFX2_11/Y OR2X2_6/gnd NAND3X1_23/A DFFSR_53/S NAND3X1
XFILL_22_DFFSR_255 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_4_NAND3X1_27 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_41_DFFSR_50 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_2_INVX1_84 INVX1_39/gnd DFFSR_34/S FILL
XFILL_3_NOR2X1_27 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_30_DFFSR_90 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_12_DFFSR_258 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_13_DFFPOSX1_26 AND2X2_38/B DFFSR_23/S FILL
XFILL_4_OAI22X1_12 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_3_NAND3X1_30 BUFX2_79/A DFFSR_6/S FILL
XDFFSR_148 INVX1_87/A CLKBUF1_31/Y BUFX2_60/Y DFFSR_175/S INVX1_88/A INVX1_67/gnd
+ DFFSR_175/S DFFSR
XFILL_2_NAND2X1_103 AND2X2_38/B DFFSR_23/S FILL
XFILL_3_OAI22X1_15 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_2_NAND3X1_33 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_14_DFFSR_40 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_4_DFFSR_145 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_1_BUFX2_75 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_1_NAND3X1_36 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_2_OAI22X1_18 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_45_DFFSR_176 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_0_NAND3X1_39 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_1_OAI22X1_21 BUFX2_98/A DFFSR_32/S FILL
XFILL_8_DFFSR_252 AND2X2_38/B DFFSR_23/S FILL
XFILL_35_DFFSR_179 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_23_DFFPOSX1_15 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_0_OAI22X1_24 BUFX2_98/A DFFSR_32/S FILL
XFILL_45_DFFSR_7 BUFX2_79/A DFFSR_7/S FILL
XFILL_25_DFFSR_182 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_49_DFFSR_57 BUFX2_79/A DFFSR_6/S FILL
XFILL_38_DFFSR_97 INVX1_1/gnd DFFSR_97/S FILL
XFILL_15_DFFSR_185 INVX1_39/gnd DFFSR_54/S FILL
XFILL_7_NAND3X1_218 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_3_DFFPOSX1_37 BUFX2_72/gnd DFFSR_201/S FILL
XINVX1_41 DFFSR_78/Q DFFSR_4/gnd INVX1_41/Y DFFSR_98/S INVX1
XDFFSR_94 DFFSR_94/Q CLKBUF1_38/Y DFFSR_15/R DFFSR_98/S DFFSR_86/Q BUFX2_77/gnd DFFSR_98/S
+ DFFSR
XFILL_22_DFFSR_47 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_5_DFFSR_54 INVX1_39/gnd DFFSR_54/S FILL
XFILL_11_DFFSR_87 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_0_NOR2X1_64 AND2X2_38/B DFFSR_59/S FILL
XFILL_48_DFFSR_103 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_38_DFFSR_106 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_8_NAND3X1_152 DFFSR_34/gnd DFFSR_1/S FILL
XINVX1_159 INVX1_159/A INVX1_3/gnd INVX1_159/Y DFFSR_79/S INVX1
XFILL_0_INVX1_9 BUFX2_99/A DFFSR_7/S FILL
XFILL_1_DFFSR_182 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_28_DFFSR_109 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_1_NAND2X1_133 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_42_DFFSR_213 INVX1_3/gnd DFFSR_23/S FILL
XFILL_4_INVX1_156 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_7_AND2X2_23 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_18_DFFSR_112 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_28_4_0 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_32_DFFSR_216 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_1_NAND2X1_3 BUFX2_99/A DFFSR_7/S FILL
XFILL_22_DFFSR_219 INVX1_67/gnd DFFSR_175/S FILL
XFILL_2_INVX1_48 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_41_DFFSR_14 INVX1_1/gnd DFFSR_53/S FILL
XFILL_19_DFFSR_94 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_30_DFFSR_54 INVX1_39/gnd DFFSR_54/S FILL
XFILL_26_6_1 INVX1_3/gnd DFFSR_23/S FILL
XFILL_12_DFFSR_222 BUFX2_72/gnd DFFSR_201/S FILL
XDFFSR_112 DFFSR_120/D DFFSR_57/CLK DFFSR_3/R DFFSR_32/S DFFSR_112/D OR2X2_4/gnd DFFSR_32/S
+ DFFSR
XFILL_22_DFFPOSX1_45 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_8_5_0 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_4_DFFSR_109 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_1_BUFX2_39 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_6_NAND3X1_248 INVX1_3/gnd DFFSR_79/S FILL
XFILL_1_OAI22X1_2 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_45_DFFSR_140 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_8_DFFSR_216 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_35_DFFSR_143 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_11_DFFSR_5 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_49_DFFSR_247 BUFX2_99/A DFFSR_7/S FILL
XFILL_25_DFFSR_146 BUFX2_79/A DFFSR_7/S FILL
XFILL_39_DFFSR_250 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_38_DFFSR_61 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_49_DFFSR_21 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_1_INVX1_193 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_15_DFFSR_149 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_7_NAND3X1_182 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_29_DFFSR_253 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_0_NAND2X1_163 INVX1_67/gnd DFFSR_201/S FILL
XDFFSR_58 DFFSR_58/Q DFFSR_8/CLK DFFSR_2/R DFFSR_3/S DFFSR_42/Q DFFSR_28/gnd DFFSR_3/S
+ DFFSR
XFILL_19_DFFSR_256 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_5_DFFSR_18 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_22_DFFSR_11 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_11_DFFSR_51 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_0_NOR2X1_28 BUFX2_98/A DFFSR_6/S FILL
XFILL_8_NAND3X1_116 DFFSR_46/gnd DFFSR_54/S FILL
XINVX1_123 BUFX2_38/Y DFFSR_34/gnd INVX1_123/Y DFFSR_1/S INVX1
XFILL_1_DFFSR_146 BUFX2_79/A DFFSR_7/S FILL
XFILL_12_DFFPOSX1_20 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_32_DFFSR_1 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_42_DFFSR_177 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_4_INVX1_120 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_46_DFFSR_68 BUFX2_98/A DFFSR_6/S FILL
XFILL_5_DFFSR_253 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_32_DFFSR_180 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_36_1_1 BUFX2_99/A DFFSR_92/S FILL
XFILL_22_DFFSR_183 INVX1_67/gnd DFFSR_175/S FILL
XFILL_2_INVX1_12 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_2_DFFSR_65 BUFX2_79/A DFFSR_7/S FILL
XFILL_19_DFFSR_58 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_30_DFFSR_18 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_12_DFFSR_186 BUFX2_99/A DFFSR_92/S FILL
XFILL_6_BUFX2_93 AND2X2_38/B DFFSR_59/S FILL
XFILL_34_3_2 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_6_NAND3X1_212 INVX1_39/gnd DFFSR_54/S FILL
XFILL_45_DFFSR_104 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_2_DFFPOSX1_31 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_8_DFFSR_180 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_35_DFFSR_107 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_49_DFFSR_211 BUFX2_7/gnd DFFSR_216/S FILL
XAND2X2_27 AOI21X1_2/Y AND2X2_27/B DFFSR_62/gnd AND2X2_27/Y DFFSR_62/S AND2X2
XFILL_25_DFFSR_110 OR2X2_3/gnd DFFSR_4/S FILL
XNAND3X1_248 XOR2X1_10/Y XOR2X1_12/B AOI21X1_64/A INVX1_3/gnd AOI21X1_68/A DFFSR_79/S
+ NAND3X1
XFILL_39_DFFSR_214 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_1_INVX1_157 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_38_DFFSR_25 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_27_DFFSR_65 BUFX2_79/A DFFSR_7/S FILL
XFILL_4_AND2X2_24 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_15_DFFSR_113 BUFX2_99/A DFFSR_92/S FILL
XFILL_7_NAND3X1_146 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_29_DFFSR_217 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_11_DFFPOSX1_50 INVX1_1/gnd DFFSR_53/S FILL
XFILL_19_DFFSR_220 BUFX2_7/gnd DFFSR_151/S FILL
XDFFSR_22 DFFSR_38/D DFFSR_92/CLK DFFSR_2/R DFFSR_32/S DFFSR_30/Q OR2X2_4/gnd DFFSR_32/S
+ DFFSR
XFILL_0_NAND2X1_127 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_11_DFFSR_15 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_1_DFFSR_110 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_21_DFFPOSX1_39 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_42_DFFSR_141 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_46_DFFSR_32 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_35_DFFSR_72 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_5_DFFSR_217 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_32_DFFSR_144 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_46_DFFSR_248 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_5_NAND3X1_242 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_22_DFFSR_147 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_2_DFFSR_29 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_36_DFFSR_251 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_19_DFFSR_22 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_6_BUFX2_57 AND2X2_38/B DFFSR_23/S FILL
XFILL_12_DFFSR_150 AND2X2_38/B DFFSR_23/S FILL
XFILL_26_DFFSR_254 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_16_DFFSR_257 INVX1_39/gnd DFFSR_34/S FILL
XFILL_20_CLKBUF1_12 AND2X2_38/B DFFSR_23/S FILL
XFILL_6_NAND3X1_176 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_43_DFFSR_79 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_19_CLKBUF1_15 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_8_DFFSR_144 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_49_DFFSR_175 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_18_CLKBUF1_18 OR2X2_1/gnd DFFSR_51/S FILL
XNAND3X1_212 NAND3X1_215/A NAND3X1_215/B AOI21X1_33/Y INVX1_39/gnd NAND3X1_218/B DFFSR_54/S
+ NAND3X1
XFILL_17_CLKBUF1_21 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_39_DFFSR_178 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_27_DFFSR_29 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_1_INVX1_121 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_16_DFFSR_69 BUFX2_98/A DFFSR_32/S FILL
XFILL_7_NAND3X1_110 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_2_DFFSR_254 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_16_CLKBUF1_24 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_29_DFFSR_181 INVX1_3/gnd DFFSR_79/S FILL
XFILL_11_DFFPOSX1_14 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_15_CLKBUF1_27 INVX1_1/gnd DFFSR_97/S FILL
XFILL_19_DFFSR_184 OR2X2_1/gnd DFFSR_51/S FILL
XNOR2X1_66 XOR2X1_1/B NOR2X1_66/B DFFSR_46/gnd NOR2X1_66/Y DFFSR_62/S NOR2X1
XFILL_14_CLKBUF1_30 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_3_XOR2X1_6 BUFX2_99/A DFFSR_7/S FILL
XFILL_23_DFFSR_8 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_51_DFFSR_86 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_13_CLKBUF1_33 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_4_NOR2X1_63 INVX1_3/gnd DFFSR_23/S FILL
XFILL_12_CLKBUF1_36 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_42_DFFSR_105 INVX1_1/gnd DFFSR_53/S FILL
XFILL_7_DFFSR_83 INVX1_3/gnd DFFSR_79/S FILL
XFILL_35_DFFSR_36 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_24_DFFSR_76 BUFX2_79/A DFFSR_7/S FILL
XFILL_11_CLKBUF1_39 INVX1_1/gnd DFFSR_53/S FILL
XFILL_5_DFFSR_181 INVX1_3/gnd DFFSR_79/S FILL
XFILL_32_DFFSR_108 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_46_DFFSR_212 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_10_CLKBUF1_42 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_5_NAND3X1_206 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_7_BUFX2_9 AND2X2_38/B DFFSR_59/S FILL
XFILL_22_DFFSR_111 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_36_DFFSR_215 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_1_DFFPOSX1_25 BUFX2_79/A DFFSR_6/S FILL
XFILL_1_AND2X2_25 INVX1_39/gnd DFFSR_54/S FILL
XFILL_6_BUFX2_21 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_5_NAND2X1_2 BUFX2_99/A DFFSR_7/S FILL
XFILL_12_DFFSR_114 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_26_DFFSR_218 BUFX2_98/A DFFSR_32/S FILL
XFILL_9_CLKBUF1_45 BUFX2_79/A DFFSR_7/S FILL
XFILL_8_CLKBUF1_48 INVX1_3/gnd DFFSR_79/S FILL
XFILL_16_DFFSR_221 AND2X2_38/B DFFSR_59/S FILL
XFILL_44_DFFSR_4 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_6_NAND3X1_140 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_10_DFFPOSX1_44 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_43_DFFSR_43 BUFX2_98/A DFFSR_6/S FILL
XFILL_32_DFFSR_83 INVX1_3/gnd DFFSR_79/S FILL
XFILL_8_DFFSR_108 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_5_OAI22X1_1 INVX1_1/gnd DFFSR_53/S FILL
XFILL_35_4_0 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_49_DFFSR_139 DFFSR_34/gnd DFFSR_34/S FILL
XNAND3X1_176 INVX1_160/A NAND3X1_176/B NAND3X1_176/C NOR3X1_6/gnd AOI21X1_28/B DFFSR_79/S
+ NAND3X1
XFILL_39_DFFSR_142 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_16_DFFSR_33 BUFX2_98/A DFFSR_32/S FILL
XFILL_22_4 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_2_DFFSR_218 BUFX2_98/A DFFSR_32/S FILL
XFILL_29_DFFSR_145 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_3_BUFX2_68 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_33_6_1 INVX1_1/gnd DFFSR_53/S FILL
XFILL_43_DFFSR_249 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_20_DFFPOSX1_33 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_19_DFFSR_148 INVX1_67/gnd DFFSR_175/S FILL
XFILL_33_DFFSR_252 AND2X2_38/B DFFSR_23/S FILL
XNOR2X1_30 NOR3X1_4/B INVX1_63/Y INVX1_3/gnd NOR2X1_30/Y DFFSR_23/S NOR2X1
XFILL_4_NAND3X1_236 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_23_DFFSR_255 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_40_DFFSR_90 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_4_NOR2X1_27 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_13_DFFSR_258 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_7_DFFSR_47 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_24_DFFSR_40 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_13_DFFSR_80 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_5_DFFSR_145 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_46_DFFSR_176 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_5_NAND3X1_170 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_9_DFFSR_252 AND2X2_38/B DFFSR_23/S FILL
XFILL_36_DFFSR_179 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_26_DFFSR_182 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_48_DFFSR_97 INVX1_1/gnd DFFSR_97/S FILL
XFILL_10_DFFSR_2 BUFX2_79/A DFFSR_7/S FILL
XFILL_8_CLKBUF1_12 AND2X2_38/B DFFSR_23/S FILL
XFILL_16_DFFSR_185 INVX1_39/gnd DFFSR_54/S FILL
XFILL_6_NAND3X1_104 AND2X2_38/B DFFSR_23/S FILL
XFILL_9_AND2X2_6 BUFX2_99/A DFFSR_7/S FILL
XFILL_7_CLKBUF1_15 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_32_DFFSR_47 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_4_DFFSR_94 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_21_DFFSR_87 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_1_NOR2X1_64 AND2X2_38/B DFFSR_59/S FILL
XFILL_6_CLKBUF1_18 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_49_DFFSR_103 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_5_CLKBUF1_21 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_43_1_1 OR2X2_4/gnd DFFSR_3/S FILL
XNAND3X1_140 AOI21X1_8/B AOI21X1_8/A OAI21X1_30/C DFFSR_1/gnd NAND2X1_64/A DFFSR_1/S
+ NAND3X1
XFILL_39_DFFSR_106 XOR2X1_4/gnd DFFSR_91/S FILL
XCLKBUF1_18 BUFX2_3/Y OR2X2_1/gnd CLKBUF1_18/Y DFFSR_51/S CLKBUF1
XFILL_5_8 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_4_CLKBUF1_24 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_2_DFFSR_182 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_29_DFFSR_109 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_3_BUFX2_32 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_43_DFFSR_213 INVX1_3/gnd DFFSR_23/S FILL
XFILL_3_CLKBUF1_27 INVX1_1/gnd DFFSR_97/S FILL
XFILL_41_3_2 BUFX2_98/A DFFSR_32/S FILL
XFILL_8_AND2X2_23 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_19_DFFSR_112 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_33_DFFSR_216 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_2_CLKBUF1_30 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_2_NAND2X1_3 BUFX2_99/A DFFSR_7/S FILL
XFILL_23_DFFSR_219 INVX1_67/gnd DFFSR_175/S FILL
XFILL_4_NAND3X1_200 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_1_CLKBUF1_33 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_51_DFFSR_14 INVX1_1/gnd DFFSR_53/S FILL
XFILL_1_INVX1_88 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_29_DFFSR_94 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_40_DFFSR_54 INVX1_39/gnd DFFSR_54/S FILL
XFILL_13_DFFSR_222 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_0_DFFPOSX1_19 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_0_CLKBUF1_36 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_7_DFFSR_11 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_13_DFFSR_44 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_5_DFFSR_109 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_0_BUFX2_79 BUFX2_79/A DFFSR_7/S FILL
XFILL_2_OAI22X1_2 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_5_NAND3X1_134 INVX1_39/gnd DFFSR_54/S FILL
XFILL_46_DFFSR_140 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_9_DFFSR_216 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_36_DFFSR_143 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_50_DFFSR_247 BUFX2_99/A DFFSR_7/S FILL
XFILL_26_DFFSR_146 BUFX2_79/A DFFSR_7/S FILL
XFILL_48_DFFSR_61 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_40_DFFSR_250 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_2_INVX1_193 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_16_DFFSR_149 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_44_4 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_30_DFFSR_253 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_20_DFFSR_256 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_4_DFFSR_58 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_32_DFFSR_11 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_10_DFFSR_91 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_21_DFFSR_51 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_19_DFFPOSX1_27 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_1_NOR2X1_28 BUFX2_98/A DFFSR_6/S FILL
XFILL_10_DFFSR_259 BUFX2_79/A DFFSR_6/S FILL
XNAND3X1_104 NOR2X1_47/Y NOR2X1_48/Y NOR2X1_49/Y AND2X2_38/B INVX1_217/A DFFSR_23/S
+ NAND3X1
XFILL_3_NAND3X1_230 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_2_DFFSR_146 BUFX2_79/A DFFSR_7/S FILL
XFILL_43_DFFSR_177 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_6_DFFSR_253 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_33_DFFSR_180 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_23_DFFSR_183 INVX1_67/gnd DFFSR_175/S FILL
XFILL_4_NAND3X1_164 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_29_DFFSR_58 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_1_INVX1_52 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_18_DFFSR_98 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_40_DFFSR_18 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_13_DFFSR_186 BUFX2_99/A DFFSR_92/S FILL
XFILL_9_DFFPOSX1_38 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_0_BUFX2_43 AND2X2_38/B DFFSR_23/S FILL
XFILL_46_DFFSR_104 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_9_DFFSR_180 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_36_DFFSR_107 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_50_DFFSR_211 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_26_DFFSR_110 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_40_DFFSR_214 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_2_INVX1_157 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_48_DFFSR_25 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_37_DFFSR_65 BUFX2_79/A DFFSR_7/S FILL
XFILL_5_AND2X2_24 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_16_DFFSR_113 BUFX2_99/A DFFSR_92/S FILL
XFILL_30_DFFSR_217 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_15_1_2 INVX1_39/gnd DFFSR_34/S FILL
XFILL_20_DFFSR_220 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_4_DFFSR_22 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_21_DFFSR_15 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_10_DFFSR_55 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_5_OAI21X1_116 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_10_DFFSR_223 INVX1_39/gnd DFFSR_34/S FILL
XFILL_3_NAND3X1_194 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_2_DFFSR_110 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_3_NOR2X1_3 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_22_DFFSR_5 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_43_DFFSR_141 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_45_DFFSR_72 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_6_DFFSR_217 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_33_DFFSR_144 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_47_DFFSR_248 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_4_NAND3X1_128 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_23_DFFSR_147 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_37_DFFSR_251 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_29_DFFSR_22 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_1_DFFSR_69 BUFX2_98/A DFFSR_32/S FILL
XFILL_1_INVX1_16 BUFX2_99/A DFFSR_7/S FILL
XFILL_18_DFFSR_62 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_13_DFFSR_150 AND2X2_38/B DFFSR_23/S FILL
XFILL_5_BUFX2_97 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_6_BUFX2_6 BUFX2_79/A DFFSR_6/S FILL
XFILL_27_DFFSR_254 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_6_NAND2X1_164 INVX1_67/gnd DFFSR_175/S FILL
XFILL_42_4_0 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_49_9 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_17_DFFSR_257 INVX1_39/gnd DFFSR_34/S FILL
XFILL_40_6_1 BUFX2_98/A DFFSR_6/S FILL
XFILL_43_DFFSR_1 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_9_DFFSR_144 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_50_DFFSR_175 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_18_DFFPOSX1_21 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_19_DFFPOSX1_3 INVX1_39/gnd DFFSR_34/S FILL
XFILL_40_DFFSR_178 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_37_DFFSR_29 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_9_DFFSR_76 BUFX2_79/A DFFSR_7/S FILL
XFILL_2_INVX1_121 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_26_DFFSR_69 BUFX2_98/A DFFSR_32/S FILL
XFILL_18_DFFPOSX1_6 AND2X2_38/B DFFSR_23/S FILL
XFILL_3_DFFSR_254 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_2_NAND3X1_224 INVX1_39/gnd DFFSR_54/S FILL
XFILL_30_DFFSR_181 INVX1_3/gnd DFFSR_79/S FILL
XFILL_17_DFFPOSX1_9 INVX1_67/gnd DFFSR_201/S FILL
XFILL_20_DFFSR_184 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_10_DFFSR_19 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_10_DFFSR_187 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_5_NOR2X1_63 INVX1_3/gnd DFFSR_23/S FILL
XFILL_3_NAND3X1_158 AND2X2_38/B DFFSR_59/S FILL
XFILL_8_DFFPOSX1_32 INVX1_67/gnd DFFSR_201/S FILL
XFILL_43_DFFSR_105 INVX1_1/gnd DFFSR_53/S FILL
XFILL_45_DFFSR_36 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_34_DFFSR_76 BUFX2_79/A DFFSR_7/S FILL
XFILL_6_DFFSR_181 INVX1_3/gnd DFFSR_79/S FILL
XFILL_33_DFFSR_108 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_47_DFFSR_212 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_23_DFFSR_111 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_1_DFFSR_33 BUFX2_98/A DFFSR_32/S FILL
XFILL_18_DFFSR_26 BUFX2_79/A DFFSR_6/S FILL
XFILL_37_DFFSR_215 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_2_AND2X2_25 INVX1_39/gnd DFFSR_54/S FILL
XFILL_13_DFFSR_114 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_6_NAND2X1_2 BUFX2_99/A DFFSR_7/S FILL
XFILL_5_BUFX2_61 AND2X2_38/B DFFSR_59/S FILL
XFILL_27_DFFSR_218 BUFX2_98/A DFFSR_32/S FILL
XFILL_10_OAI22X1_7 AND2X2_38/B DFFSR_59/S FILL
XFILL_6_NAND2X1_128 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_17_DFFSR_221 AND2X2_38/B DFFSR_59/S FILL
XFILL_50_1_1 DFFSR_4/gnd DFFSR_4/S FILL
XXOR2X1_3 XOR2X1_3/A XOR2X1_3/B OR2X2_2/gnd XOR2X1_3/Y DFFSR_216/S XOR2X1
XFILL_9_AOI21X1_53 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_9_DFFSR_108 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_42_DFFSR_83 INVX1_3/gnd DFFSR_79/S FILL
XNAND2X1_164 NAND2X1_163/B INVX1_208/Y INVX1_67/gnd AOI21X1_58/A DFFSR_175/S NAND2X1
XFILL_48_3_2 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_6_OAI22X1_1 INVX1_1/gnd DFFSR_53/S FILL
XFILL_4_OAI21X1_110 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_50_DFFSR_139 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_8_AOI21X1_56 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_27_DFFPOSX1_40 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_40_DFFSR_142 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_9_DFFSR_40 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_26_1 AND2X2_38/B DFFSR_23/S FILL
XFILL_26_DFFSR_33 BUFX2_98/A DFFSR_32/S FILL
XFILL_7_AOI21X1_59 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_15_DFFSR_73 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_2_NAND3X1_188 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_3_DFFSR_218 BUFX2_98/A DFFSR_32/S FILL
XFILL_30_DFFSR_145 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_6_AOI21X1_62 INVX1_3/gnd DFFSR_23/S FILL
XFILL_44_DFFSR_249 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_20_DFFSR_148 INVX1_67/gnd DFFSR_175/S FILL
XFILL_5_AOI21X1_65 INVX1_3/gnd DFFSR_23/S FILL
XFILL_34_DFFSR_252 AND2X2_38/B DFFSR_23/S FILL
XFILL_10_DFFSR_151 XOR2X1_1/gnd DFFSR_151/S FILL
XAOI21X1_62 BUFX2_7/Y OR2X2_1/A NOR3X1_1/A INVX1_3/gnd NOR2X1_76/A DFFSR_23/S AOI21X1
XFILL_4_AOI21X1_68 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_24_DFFSR_255 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_50_DFFSR_90 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_5_NOR2X1_27 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_3_NAND3X1_122 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_14_DFFSR_258 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_3_AOI21X1_71 BUFX2_99/A DFFSR_92/S FILL
XFILL_16_2_0 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_34_DFFSR_40 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_23_DFFSR_80 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_6_DFFSR_87 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_5_NAND2X1_158 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_6_DFFSR_145 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_14_4_1 INVX1_39/gnd DFFSR_54/S FILL
XFILL_47_DFFSR_176 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_37_DFFSR_179 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_8_OR2X2_4 OR2X2_4/gnd DFFSR_32/S FILL
XBUFX2_65 BUFX2_60/A DFFSR_8/gnd BUFX2_65/Y DFFSR_60/S BUFX2
XFILL_0_DFFSR_255 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_5_BUFX2_25 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_17_DFFPOSX1_15 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_12_6_2 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_27_DFFSR_182 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_17_DFFSR_185 INVX1_39/gnd DFFSR_54/S FILL
XFILL_34_DFFSR_8 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_15_NOR3X1_4 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_1_NAND3X1_218 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_3_INVX1_81 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_9_AOI21X1_17 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_31_DFFSR_87 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_42_DFFSR_47 BUFX2_77/gnd DFFSR_98/S FILL
XNAND2X1_128 BUFX2_53/Y INVX1_154/A BUFX2_72/gnd OAI21X1_97/C DFFSR_276/S NAND2X1
XFILL_2_NOR2X1_64 AND2X2_38/B DFFSR_59/S FILL
XFILL_50_DFFSR_103 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_8_AOI21X1_20 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_7_DFFPOSX1_3 INVX1_39/gnd DFFSR_34/S FILL
XFILL_40_DFFSR_106 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_6_DFFPOSX1_6 AND2X2_38/B DFFSR_23/S FILL
XFILL_7_AOI21X1_23 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_9_5 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_15_DFFSR_37 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_2_NAND3X1_152 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_3_DFFSR_182 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_2_BUFX2_72 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_5_DFFPOSX1_9 INVX1_67/gnd DFFSR_201/S FILL
XFILL_30_DFFSR_109 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_44_DFFSR_213 INVX1_3/gnd DFFSR_23/S FILL
XFILL_6_AOI21X1_26 DFFSR_62/gnd DFFSR_208/S FILL
XDFFPOSX1_6 NOR3X1_4/B CLKBUF1_43/Y NAND2X1_54/Y AND2X2_38/B DFFSR_23/S DFFPOSX1
XFILL_9_AND2X2_23 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_20_DFFSR_112 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_7_DFFPOSX1_26 AND2X2_38/B DFFSR_23/S FILL
XFILL_5_AOI21X1_29 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_34_DFFSR_216 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_10_DFFSR_115 INVX1_1/gnd DFFSR_97/S FILL
XAOI21X1_26 AOI21X1_26/A AOI21X1_26/B AOI21X1_26/C DFFSR_62/gnd AOI21X1_26/Y DFFSR_208/S
+ AOI21X1
XFILL_3_NAND2X1_3 BUFX2_99/A DFFSR_7/S FILL
XFILL_4_AOI21X1_32 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_24_DFFSR_219 INVX1_67/gnd DFFSR_175/S FILL
XFILL_39_DFFSR_94 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_50_DFFSR_54 INVX1_39/gnd DFFSR_54/S FILL
XFILL_14_DFFSR_222 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_3_AOI21X1_35 INVX1_39/gnd DFFSR_54/S FILL
XFILL_2_AOI21X1_38 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_16_DFFPOSX1_45 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_0_AND2X2_3 INVX1_1/gnd DFFSR_53/S FILL
XFILL_5_NAND2X1_122 INVX1_67/gnd DFFSR_175/S FILL
XFILL_23_DFFSR_44 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_6_DFFSR_51 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_6_DFFSR_109 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_12_DFFSR_84 BUFX2_99/A DFFSR_7/S FILL
XFILL_1_AOI21X1_41 INVX1_39/gnd DFFSR_34/S FILL
XFILL_3_OAI22X1_2 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_0_NAND3X1_248 INVX1_3/gnd DFFSR_79/S FILL
XFILL_47_DFFSR_140 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_0_AOI21X1_44 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_22_1_2 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_37_DFFSR_143 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_0_DFFSR_219 INVX1_67/gnd DFFSR_175/S FILL
XBUFX2_29 BUFX2_27/A BUFX2_8/gnd BUFX2_29/Y DFFSR_51/S BUFX2
XFILL_4_0_1 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_3_OAI21X1_104 INVX1_67/gnd DFFSR_201/S FILL
XFILL_27_DFFSR_146 BUFX2_79/A DFFSR_7/S FILL
XFILL_31_6 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_26_DFFPOSX1_34 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_41_DFFSR_250 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_3_INVX1_193 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_17_DFFSR_149 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_48_1 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_8_OAI21X1_68 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_1_NAND3X1_182 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_31_DFFSR_253 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_2_2_2 INVX1_67/gnd DFFSR_201/S FILL
XFILL_21_DFFSR_256 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_7_OAI21X1_71 INVX1_3/gnd DFFSR_79/S FILL
XFILL_6_NAND2X1_89 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_3_INVX1_45 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_42_DFFSR_11 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_3_DFFSR_98 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_20_DFFSR_91 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_31_DFFSR_51 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_2_NOR2X1_28 BUFX2_98/A DFFSR_6/S FILL
XFILL_5_NAND2X1_92 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_6_OAI21X1_74 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_11_DFFSR_259 BUFX2_79/A DFFSR_6/S FILL
XNAND2X1_89 AOI22X1_24/A AOI22X1_24/B DFFSR_46/gnd AOI21X1_22/C DFFSR_54/S NAND2X1
XFILL_5_OAI21X1_77 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_4_NAND2X1_95 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_2_NAND3X1_116 DFFSR_46/gnd DFFSR_54/S FILL
XOAI21X1_74 OAI21X1_74/A AOI21X1_23/Y INVX1_163/A DFFSR_46/gnd OAI21X1_74/Y DFFSR_62/S
+ OAI21X1
XFILL_3_DFFSR_146 BUFX2_79/A DFFSR_7/S FILL
XFILL_3_NAND2X1_98 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_2_BUFX2_36 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_4_OAI21X1_80 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_44_DFFSR_177 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_3_OAI21X1_83 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_7_DFFSR_253 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_49_4_0 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_4_NAND2X1_152 INVX1_1/gnd DFFSR_97/S FILL
XFILL_34_DFFSR_180 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_2_OAI21X1_86 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_21_DFFSR_2 BUFX2_79/A DFFSR_7/S FILL
XFILL_24_DFFSR_183 INVX1_67/gnd DFFSR_175/S FILL
XFILL_1_OAI21X1_89 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_39_DFFSR_58 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_50_DFFSR_18 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_0_INVX1_92 AND2X2_38/B DFFSR_23/S FILL
XFILL_28_DFFSR_98 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_47_6_1 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_14_DFFSR_186 BUFX2_99/A DFFSR_92/S FILL
XFILL_0_OAI21X1_92 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_6_DFFSR_15 OR2X2_3/gnd DFFSR_4/S FILL
XBUFX2_7 BUFX2_7/A BUFX2_7/gnd BUFX2_7/Y DFFSR_151/S BUFX2
XFILL_12_DFFSR_48 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_5_BUFX2_3 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_47_DFFSR_104 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_0_NAND3X1_212 INVX1_39/gnd DFFSR_54/S FILL
XFILL_37_DFFSR_107 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_51_DFFSR_211 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_0_DFFSR_183 INVX1_67/gnd DFFSR_175/S FILL
XFILL_27_DFFSR_110 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_41_DFFSR_214 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_3_INVX1_157 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_47_DFFSR_65 BUFX2_79/A DFFSR_7/S FILL
XFILL_6_AND2X2_24 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_17_DFFSR_113 BUFX2_99/A DFFSR_92/S FILL
XFILL_8_OAI21X1_32 AND2X2_38/B DFFSR_59/S FILL
XFILL_31_DFFSR_217 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_1_NAND3X1_146 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_0_NAND2X1_4 BUFX2_98/A DFFSR_6/S FILL
XFILL_7_OAI21X1_35 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_21_DFFSR_220 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_6_NAND2X1_53 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_31_DFFSR_15 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_20_DFFSR_55 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_3_DFFSR_62 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_6_DFFPOSX1_20 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_3_NAND2X1_182 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_5_NAND2X1_56 AND2X2_38/B DFFSR_59/S FILL
XFILL_6_OAI21X1_38 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_11_DFFSR_223 INVX1_39/gnd DFFSR_34/S FILL
XNAND2X1_53 AOI21X1_1/A AOI21X1_1/B DFFSR_62/gnd AOI21X1_2/A DFFSR_62/S NAND2X1
XFILL_5_OAI21X1_41 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_4_NAND2X1_59 DFFSR_62/gnd DFFSR_208/S FILL
XOAI21X1_38 INVX1_144/A AOI22X1_18/Y OAI21X1_38/C OR2X2_1/gnd AOI21X1_11/C DFFSR_59/S
+ OAI21X1
XFILL_3_DFFSR_110 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_3_NAND2X1_62 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_4_OAI21X1_44 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_0_OAI22X1_3 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_44_DFFSR_141 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_15_DFFPOSX1_39 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_2_NAND2X1_65 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_3_OAI21X1_47 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_7_DFFSR_217 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_4_NAND2X1_116 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_34_DFFSR_144 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_2_OAI21X1_50 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_1_NAND2X1_68 AND2X2_38/B DFFSR_23/S FILL
XFILL_48_DFFSR_248 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_24_DFFSR_147 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_0_NAND2X1_71 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_1_OAI21X1_53 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_0_INVX1_194 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_38_DFFSR_251 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_39_DFFSR_22 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_0_INVX1_56 BUFX2_98/A DFFSR_6/S FILL
XFILL_10_AOI22X1_19 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_28_DFFSR_62 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_14_DFFSR_150 AND2X2_38/B DFFSR_23/S FILL
XFILL_28_DFFSR_254 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_0_OAI21X1_56 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_25_DFFPOSX1_28 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_18_DFFSR_257 INVX1_39/gnd DFFSR_34/S FILL
XFILL_9_AOI22X1_22 INVX1_3/gnd DFFSR_79/S FILL
XFILL_12_DFFSR_12 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_8_AOI22X1_25 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_0_NAND3X1_176 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_7_AOI22X1_28 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_5_DFFPOSX1_50 INVX1_1/gnd DFFSR_53/S FILL
XFILL_0_DFFSR_147 DFFSR_1/gnd DFFSR_1/S FILL
XDFFSR_257 DFFSR_1/D DFFSR_1/CLK DFFSR_257/R DFFSR_34/S DFFSR_257/D INVX1_39/gnd DFFSR_34/S
+ DFFSR
XFILL_41_DFFSR_178 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_3_INVX1_121 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_47_DFFSR_29 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_36_DFFSR_69 BUFX2_98/A DFFSR_32/S FILL
XFILL_4_DFFSR_254 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_1_NAND3X1_110 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_31_DFFSR_181 INVX1_3/gnd DFFSR_79/S FILL
XFILL_23_2_0 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_6_NAND2X1_17 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_21_DFFSR_184 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_3_DFFSR_26 BUFX2_79/A DFFSR_6/S FILL
XFILL_20_DFFSR_19 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_3_NAND2X1_146 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_5_NAND2X1_20 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_11_DFFSR_187 DFFSR_1/gnd DFFSR_81/S FILL
XNAND2X1_17 DFFSR_116/D NOR2X1_5/Y OR2X2_6/gnd OAI21X1_4/C DFFSR_92/S NAND2X1
XFILL_4_NAND2X1_23 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_21_4_1 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_6_NOR2X1_63 INVX1_3/gnd DFFSR_23/S FILL
XFILL_3_NAND2X1_26 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_2_NOR2X1_7 BUFX2_98/A DFFSR_32/S FILL
XFILL_3_3_0 INVX1_67/gnd DFFSR_175/S FILL
XFILL_9_DFFSR_1 DFFSR_1/gnd DFFSR_1/S FILL
XDFFPOSX1_20 INVX1_169/A CLKBUF1_47/Y OAI22X1_51/Y DFFSR_46/gnd DFFSR_62/S DFFPOSX1
XFILL_12_DFFSR_9 BUFX2_79/A DFFSR_6/S FILL
XFILL_44_DFFSR_105 INVX1_1/gnd DFFSR_53/S FILL
XFILL_44_DFFSR_76 BUFX2_79/A DFFSR_7/S FILL
XFILL_2_NAND2X1_29 INVX1_3/gnd DFFSR_23/S FILL
XFILL_19_6_2 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_3_OAI21X1_11 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_7_DFFSR_181 INVX1_3/gnd DFFSR_79/S FILL
XFILL_34_DFFSR_108 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_48_DFFSR_212 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_1_NAND2X1_32 INVX1_3/gnd DFFSR_79/S FILL
XFILL_2_OAI21X1_14 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_1_5_1 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_24_DFFSR_111 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_8_NAND3X1_88 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_0_NAND2X1_35 INVX1_67/gnd DFFSR_201/S FILL
XFILL_1_OAI21X1_17 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_28_DFFSR_26 BUFX2_79/A DFFSR_6/S FILL
XFILL_0_INVX1_20 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_0_DFFSR_73 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_38_DFFSR_215 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_0_INVX1_158 INVX1_39/gnd DFFSR_34/S FILL
XFILL_17_DFFSR_66 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_3_AND2X2_25 INVX1_39/gnd DFFSR_54/S FILL
XFILL_14_DFFSR_114 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_7_NAND3X1_91 AND2X2_38/B DFFSR_59/S FILL
XFILL_28_DFFSR_218 BUFX2_98/A DFFSR_32/S FILL
XFILL_0_OAI21X1_20 AND2X2_38/B DFFSR_23/S FILL
XFILL_11_OAI22X1_7 AND2X2_38/B DFFSR_59/S FILL
XFILL_6_NAND3X1_94 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_18_DFFSR_221 AND2X2_38/B DFFSR_59/S FILL
XFILL_7_OR2X2_1 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_5_NAND3X1_97 AND2X2_38/B DFFSR_59/S FILL
XFILL_4_XOR2X1_3 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_0_NAND3X1_140 DFFSR_1/gnd DFFSR_1/S FILL
XNAND3X1_94 DFFSR_204/D BUFX2_27/Y NOR2X1_31/Y DFFSR_62/gnd NAND3X1_94/Y DFFSR_208/S
+ NAND3X1
XFILL_33_DFFSR_5 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_7_OAI22X1_1 INVX1_1/gnd DFFSR_53/S FILL
XFILL_5_DFFPOSX1_14 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_0_DFFSR_111 DFFSR_8/gnd DFFSR_8/S FILL
XDFFSR_221 DFFSR_229/D CLKBUF1_12/Y BUFX2_70/Y DFFSR_59/S INVX1_92/A AND2X2_38/B DFFSR_59/S
+ DFFSR
XFILL_2_NAND2X1_176 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_41_DFFSR_142 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_8_DFFSR_80 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_36_DFFSR_33 BUFX2_98/A DFFSR_32/S FILL
XFILL_25_DFFSR_73 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_4_DFFSR_218 BUFX2_98/A DFFSR_32/S FILL
XFILL_31_DFFSR_145 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_45_DFFSR_249 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_21_DFFSR_148 INVX1_67/gnd DFFSR_175/S FILL
XFILL_14_DFFPOSX1_33 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_35_DFFSR_252 AND2X2_38/B DFFSR_23/S FILL
XFILL_11_DFFSR_151 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_3_NAND2X1_110 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_25_DFFSR_255 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_6_NOR2X1_27 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_29_1_2 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_15_DFFSR_258 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_0_NOR3X1_4 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_1_AOI22X1_10 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_10_OAI22X1_31 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_0_AOI22X1_13 AND2X2_38/B DFFSR_23/S FILL
XFILL_44_DFFSR_40 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_7_DFFSR_145 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_33_DFFSR_80 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_24_DFFPOSX1_22 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_48_DFFSR_176 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_8_NAND3X1_52 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_9_OAI22X1_34 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_9_2_2 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_0_DFFSR_37 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_8_NAND3X1_225 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_38_DFFSR_179 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_0_INVX1_122 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_17_DFFSR_30 BUFX2_98/A DFFSR_32/S FILL
XFILL_7_NAND3X1_55 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_4_BUFX2_65 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_1_DFFSR_255 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_8_OAI22X1_37 INVX1_3/gnd DFFSR_23/S FILL
XFILL_4_DFFPOSX1_44 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_28_DFFSR_182 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_6_NAND3X1_58 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_7_OAI22X1_40 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_18_DFFSR_185 INVX1_39/gnd DFFSR_54/S FILL
XFILL_5_NAND3X1_61 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_6_OAI22X1_43 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_0_NAND3X1_104 AND2X2_38/B DFFSR_23/S FILL
XNAND3X1_58 DFFSR_8/Q NOR2X1_4/Y BUFX2_17/Y DFFSR_28/gnd AND2X2_13/B DFFSR_3/S NAND3X1
XFILL_4_NAND3X1_64 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_5_OAI22X1_46 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_41_DFFSR_87 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_3_NOR2X1_64 AND2X2_38/B DFFSR_59/S FILL
XOAI22X1_43 INVX1_104/Y OAI22X1_43/B INVX1_105/Y OAI22X1_43/D DFFSR_62/gnd NOR2X1_53/B
+ DFFSR_208/S OAI22X1
XFILL_3_NAND3X1_67 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_4_OAI22X1_49 OR2X2_1/gnd DFFSR_59/S FILL
XDFFSR_185 INVX1_61/A CLKBUF1_17/Y BUFX2_69/Y DFFSR_54/S DFFSR_169/Q INVX1_39/gnd
+ DFFSR_54/S DFFSR
XFILL_2_NAND2X1_140 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_41_DFFSR_106 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_2_NAND3X1_70 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_3_OAI22X1_52 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_25_DFFSR_37 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_8_DFFSR_44 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_14_DFFSR_77 BUFX2_98/A DFFSR_32/S FILL
XFILL_4_DFFSR_182 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_31_DFFSR_109 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_1_NAND3X1_73 INVX1_1/gnd DFFSR_97/S FILL
XFILL_54_6_1 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_45_DFFSR_213 INVX1_3/gnd DFFSR_23/S FILL
XNAND2X1_6 NOR2X1_4/Y NOR2X1_1/Y BUFX2_98/A OAI22X1_6/B DFFSR_32/S NAND2X1
XFILL_21_DFFSR_112 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_0_NAND3X1_76 INVX1_1/gnd DFFSR_53/S FILL
XFILL_35_DFFSR_216 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_0_AND2X2_26 INVX1_1/gnd DFFSR_97/S FILL
XFILL_11_DFFSR_115 INVX1_1/gnd DFFSR_97/S FILL
XFILL_4_NAND2X1_3 BUFX2_99/A DFFSR_7/S FILL
XFILL_25_DFFSR_219 INVX1_67/gnd DFFSR_175/S FILL
XFILL_0_DFFSR_8 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_49_DFFSR_94 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_15_DFFSR_222 BUFX2_72/gnd DFFSR_201/S FILL
XOAI22X1_5 INVX1_12/Y OAI22X1_2/B INVX1_13/Y OAI22X1_2/D DFFSR_4/gnd NOR2X1_9/A DFFSR_98/S
+ OAI22X1
XINVX1_78 INVX1_78/A DFFSR_46/gnd INVX1_78/Y DFFSR_62/S INVX1
XFILL_5_DFFSR_91 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_7_DFFSR_109 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_33_DFFSR_44 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_22_DFFSR_84 BUFX2_99/A DFFSR_7/S FILL
XFILL_9_NAND3X1_13 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_4_OAI22X1_2 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_48_DFFSR_140 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_8_NAND3X1_16 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_38_DFFSR_143 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_8_NAND3X1_189 BUFX2_7/gnd DFFSR_151/S FILL
XINVX1_196 INVX1_196/A DFFSR_1/gnd INVX1_196/Y DFFSR_81/S INVX1
XFILL_1_DFFSR_219 INVX1_67/gnd DFFSR_175/S FILL
XFILL_7_NAND3X1_19 BUFX2_99/A DFFSR_92/S FILL
XFILL_4_BUFX2_29 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_28_DFFSR_146 BUFX2_79/A DFFSR_7/S FILL
XFILL_1_NAND2X1_170 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_42_DFFSR_250 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_6_NAND3X1_22 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_18_DFFSR_149 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_32_DFFSR_253 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_5_NAND3X1_25 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_22_DFFSR_256 DFFSR_8/gnd DFFSR_60/S FILL
XNAND3X1_22 DFFSR_67/Q BUFX2_18/Y NOR2X1_2/Y OR2X2_6/gnd NAND3X1_22/Y DFFSR_53/S NAND3X1
XFILL_4_NAND3X1_28 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_5_OAI22X1_10 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_30_DFFSR_91 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_41_DFFSR_51 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_2_INVX1_85 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_3_NOR2X1_28 BUFX2_98/A DFFSR_6/S FILL
XFILL_13_DFFPOSX1_27 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_3_NAND3X1_31 BUFX2_79/A DFFSR_6/S FILL
XFILL_12_DFFSR_259 BUFX2_79/A DFFSR_6/S FILL
XDFFSR_149 INVX1_94/A CLKBUF1_10/Y BUFX2_62/Y DFFSR_276/S INVX1_95/A BUFX2_72/gnd
+ DFFSR_276/S DFFSR
XFILL_4_OAI22X1_13 INVX1_1/gnd DFFSR_53/S FILL
XFILL_2_NAND2X1_104 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_2_NAND3X1_34 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_3_OAI22X1_16 AND2X2_38/B DFFSR_59/S FILL
XFILL_14_DFFSR_41 BUFX2_98/A DFFSR_6/S FILL
XFILL_4_DFFSR_146 BUFX2_79/A DFFSR_7/S FILL
XFILL_1_BUFX2_76 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_2_OAI22X1_19 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_1_NAND3X1_37 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_45_DFFSR_177 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_1_OAI22X1_22 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_0_NAND3X1_40 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_8_DFFSR_253 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_35_DFFSR_180 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_23_DFFPOSX1_16 INVX1_67/gnd DFFSR_175/S FILL
XFILL_0_OAI22X1_25 INVX1_39/gnd DFFSR_54/S FILL
XFILL_25_DFFSR_183 INVX1_67/gnd DFFSR_175/S FILL
XFILL_45_DFFSR_8 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_49_DFFSR_58 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_38_DFFSR_98 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_15_DFFSR_186 BUFX2_99/A DFFSR_92/S FILL
XFILL_7_NAND3X1_219 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_3_DFFPOSX1_38 OR2X2_1/gnd DFFSR_51/S FILL
XINVX1_42 DFFSR_38/D OR2X2_4/gnd INVX1_42/Y DFFSR_32/S INVX1
XFILL_5_DFFSR_55 DFFSR_4/gnd DFFSR_4/S FILL
XDFFSR_95 DFFSR_95/Q CLKBUF1_38/Y DFFSR_15/R DFFSR_5/S INVX1_47/A DFFSR_5/gnd DFFSR_5/S
+ DFFSR
XFILL_22_DFFSR_48 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_11_DFFSR_88 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_0_NOR2X1_65 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_48_DFFSR_104 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_30_2_0 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_38_DFFSR_107 OR2X2_6/gnd DFFSR_92/S FILL
XINVX1_160 INVX1_160/A XOR2X1_4/gnd INVX1_160/Y DFFSR_97/S INVX1
XFILL_8_NAND3X1_153 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_1_DFFSR_183 INVX1_67/gnd DFFSR_175/S FILL
XFILL_28_DFFSR_110 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_1_NAND2X1_134 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_42_DFFSR_214 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_4_INVX1_157 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_7_AND2X2_24 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_18_DFFSR_113 BUFX2_99/A DFFSR_92/S FILL
XFILL_28_4_1 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_32_DFFSR_217 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_1_NAND2X1_4 BUFX2_98/A DFFSR_6/S FILL
XFILL_22_DFFSR_220 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_41_DFFSR_15 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_30_DFFSR_55 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_2_INVX1_49 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_19_DFFSR_95 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_26_6_2 INVX1_3/gnd DFFSR_23/S FILL
XFILL_12_DFFSR_223 INVX1_39/gnd DFFSR_34/S FILL
XDFFSR_113 INVX1_9/A CLKBUF1_40/Y BUFX2_49/Y DFFSR_92/S DFFSR_105/Q BUFX2_99/A DFFSR_92/S
+ DFFSR
XFILL_22_DFFPOSX1_46 INVX1_39/gnd DFFSR_34/S FILL
XFILL_8_5_1 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_4_DFFSR_110 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_6_NAND3X1_249 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_1_OAI22X1_3 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_1_BUFX2_40 INVX1_1/gnd DFFSR_97/S FILL
XFILL_45_DFFSR_141 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_8_DFFSR_217 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_35_DFFSR_144 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_49_DFFSR_248 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_11_DFFSR_6 BUFX2_79/A DFFSR_6/S FILL
XFILL_25_DFFSR_147 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_1_INVX1_194 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_39_DFFSR_251 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_49_DFFSR_22 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_38_DFFSR_62 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_15_DFFSR_150 AND2X2_38/B DFFSR_23/S FILL
XFILL_7_NAND3X1_183 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_29_DFFSR_254 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_0_NAND2X1_164 INVX1_67/gnd DFFSR_175/S FILL
XFILL_5_DFFSR_19 DFFSR_28/gnd DFFSR_8/S FILL
XDFFSR_59 DFFSR_51/D CLKBUF1_18/Y DFFSR_73/R DFFSR_59/S DFFSR_59/D AND2X2_38/B DFFSR_59/S
+ DFFSR
XFILL_19_DFFSR_257 INVX1_39/gnd DFFSR_34/S FILL
XFILL_22_DFFSR_12 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_11_DFFSR_52 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_0_NOR2X1_29 DFFSR_28/gnd DFFSR_3/S FILL
XINVX1_124 BUFX2_38/Y DFFSR_34/gnd INVX1_124/Y DFFSR_1/S INVX1
XFILL_8_NAND3X1_117 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_1_DFFSR_147 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_12_DFFPOSX1_21 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_32_DFFSR_2 BUFX2_79/A DFFSR_7/S FILL
XFILL_42_DFFSR_178 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_4_INVX1_121 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_46_DFFSR_69 BUFX2_98/A DFFSR_32/S FILL
XFILL_5_DFFSR_254 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_32_DFFSR_181 INVX1_3/gnd DFFSR_79/S FILL
XFILL_36_1_2 BUFX2_99/A DFFSR_92/S FILL
XFILL_22_DFFSR_184 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_30_DFFSR_19 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_2_INVX1_13 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_2_DFFSR_66 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_19_DFFSR_59 AND2X2_38/B DFFSR_59/S FILL
XFILL_6_BUFX2_94 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_12_DFFSR_187 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_22_DFFPOSX1_10 INVX1_67/gnd DFFSR_201/S FILL
XFILL_20_CLKBUF1_49 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_6_NAND3X1_213 INVX1_39/gnd DFFSR_54/S FILL
XFILL_45_DFFSR_105 INVX1_1/gnd DFFSR_53/S FILL
XFILL_2_DFFPOSX1_32 INVX1_67/gnd DFFSR_201/S FILL
XFILL_8_DFFSR_181 INVX1_3/gnd DFFSR_79/S FILL
XFILL_35_DFFSR_108 OR2X2_6/gnd DFFSR_92/S FILL
XAND2X2_28 BUFX2_8/Y OR2X2_1/A BUFX2_8/gnd AND2X2_28/Y DFFSR_51/S AND2X2
XFILL_49_DFFSR_212 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_25_DFFSR_111 DFFSR_8/gnd DFFSR_8/S FILL
XNAND3X1_249 AOI21X1_71/B XNOR2X1_4/Y AOI21X1_71/A OR2X2_6/gnd NAND2X1_182/B DFFSR_92/S
+ NAND3X1
XFILL_39_DFFSR_215 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_1_INVX1_158 INVX1_39/gnd DFFSR_34/S FILL
XFILL_27_DFFSR_66 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_38_DFFSR_26 BUFX2_79/A DFFSR_6/S FILL
XFILL_4_AND2X2_25 INVX1_39/gnd DFFSR_54/S FILL
XFILL_15_DFFSR_114 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_7_NAND3X1_147 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_29_DFFSR_218 BUFX2_98/A DFFSR_32/S FILL
XFILL_0_NAND2X1_128 BUFX2_72/gnd DFFSR_276/S FILL
XDFFSR_23 DFFSR_23/Q CLKBUF1_18/Y DFFSR_1/R DFFSR_23/S DFFSR_23/D AND2X2_38/B DFFSR_23/S
+ DFFSR
XFILL_19_DFFSR_221 AND2X2_38/B DFFSR_59/S FILL
XFILL_11_DFFSR_16 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_8_OAI22X1_1 INVX1_1/gnd DFFSR_53/S FILL
XFILL_1_DFFSR_111 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_21_DFFPOSX1_40 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_42_DFFSR_142 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_46_DFFSR_33 BUFX2_98/A DFFSR_32/S FILL
XFILL_35_DFFSR_73 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_5_DFFSR_218 BUFX2_98/A DFFSR_32/S FILL
XFILL_32_DFFSR_145 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_46_DFFSR_249 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_5_NAND3X1_243 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_22_DFFSR_148 INVX1_67/gnd DFFSR_175/S FILL
XFILL_2_DFFSR_30 BUFX2_98/A DFFSR_32/S FILL
XFILL_19_DFFSR_23 AND2X2_38/B DFFSR_23/S FILL
XFILL_36_DFFSR_252 AND2X2_38/B DFFSR_23/S FILL
XFILL_12_DFFSR_151 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_6_BUFX2_58 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_26_DFFSR_255 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_16_DFFSR_258 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_20_CLKBUF1_13 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_6_NAND3X1_177 AND2X2_38/B DFFSR_59/S FILL
XFILL_19_CLKBUF1_16 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_8_DFFSR_145 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_43_DFFSR_80 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_49_DFFSR_176 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_18_CLKBUF1_19 BUFX2_8/gnd DFFSR_81/S FILL
XNAND3X1_213 AOI21X1_26/Y NAND3X1_218/B XOR2X1_8/A INVX1_39/gnd NAND3X1_217/B DFFSR_54/S
+ NAND3X1
XFILL_17_CLKBUF1_22 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_39_DFFSR_179 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_1_INVX1_122 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_16_DFFSR_70 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_27_DFFSR_30 BUFX2_98/A DFFSR_32/S FILL
XFILL_7_NAND3X1_111 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_2_DFFSR_255 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_16_CLKBUF1_25 INVX1_67/gnd DFFSR_201/S FILL
XFILL_29_DFFSR_182 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_11_DFFPOSX1_15 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_15_CLKBUF1_28 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_19_DFFSR_185 INVX1_39/gnd DFFSR_54/S FILL
XNOR2X1_67 INVX1_153/A INVX1_141/Y INVX1_67/gnd NOR2X1_67/Y DFFSR_175/S NOR2X1
XFILL_14_CLKBUF1_31 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_3_XOR2X1_7 BUFX2_98/A DFFSR_6/S FILL
XFILL_13_CLKBUF1_34 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_23_DFFSR_9 BUFX2_79/A DFFSR_6/S FILL
XFILL_4_NOR2X1_64 AND2X2_38/B DFFSR_59/S FILL
XFILL_12_CLKBUF1_37 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_42_DFFSR_106 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_35_DFFSR_37 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_7_DFFSR_84 BUFX2_99/A DFFSR_7/S FILL
XFILL_24_DFFSR_77 BUFX2_98/A DFFSR_32/S FILL
XFILL_11_CLKBUF1_40 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_5_DFFSR_182 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_32_DFFSR_109 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_46_DFFSR_213 INVX1_3/gnd DFFSR_23/S FILL
XFILL_10_CLKBUF1_43 AND2X2_38/B DFFSR_23/S FILL
XFILL_5_NAND3X1_207 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_22_DFFSR_112 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_36_DFFSR_216 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_1_DFFPOSX1_26 AND2X2_38/B DFFSR_23/S FILL
XFILL_1_AND2X2_26 INVX1_1/gnd DFFSR_97/S FILL
XFILL_12_DFFSR_115 INVX1_1/gnd DFFSR_97/S FILL
XFILL_5_NAND2X1_3 BUFX2_99/A DFFSR_7/S FILL
XFILL_6_BUFX2_22 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_26_DFFSR_219 INVX1_67/gnd DFFSR_175/S FILL
XFILL_9_CLKBUF1_46 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_16_DFFSR_222 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_8_CLKBUF1_49 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_44_DFFSR_5 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_16_NOR3X1_1 INVX1_3/gnd DFFSR_79/S FILL
XFILL_37_2_0 BUFX2_99/A DFFSR_7/S FILL
XFILL_6_NAND3X1_141 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_10_DFFPOSX1_45 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_8_DFFSR_109 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_43_DFFSR_44 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_32_DFFSR_84 BUFX2_99/A DFFSR_7/S FILL
XFILL_4_INVX1_78 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_5_OAI22X1_2 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_35_4_1 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_49_DFFSR_140 DFFSR_62/gnd DFFSR_208/S FILL
XNAND3X1_177 AOI21X1_27/C AOI21X1_28/B AOI21X1_28/A AND2X2_38/B AOI21X1_21/A DFFSR_59/S
+ NAND3X1
XFILL_39_DFFSR_143 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_22_5 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_16_DFFSR_34 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_2_DFFSR_219 INVX1_67/gnd DFFSR_175/S FILL
XFILL_3_BUFX2_69 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_29_DFFSR_146 BUFX2_79/A DFFSR_7/S FILL
XFILL_33_6_2 INVX1_1/gnd DFFSR_53/S FILL
XFILL_43_DFFSR_250 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_19_DFFSR_149 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_20_DFFPOSX1_34 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_33_DFFSR_253 DFFSR_34/gnd DFFSR_1/S FILL
XNOR2X1_31 NOR3X1_3/A NOR3X1_3/B INVX1_39/gnd NOR2X1_31/Y DFFSR_54/S NOR2X1
XFILL_23_DFFSR_256 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_4_NAND3X1_237 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_40_DFFSR_91 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_51_DFFSR_51 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_4_NOR2X1_28 BUFX2_98/A DFFSR_6/S FILL
XFILL_13_DFFSR_259 BUFX2_79/A DFFSR_6/S FILL
XFILL_7_DFFSR_48 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_24_DFFSR_41 BUFX2_98/A DFFSR_6/S FILL
XFILL_5_DFFSR_146 BUFX2_79/A DFFSR_7/S FILL
XFILL_13_DFFSR_81 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_5_NAND3X1_171 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_46_DFFSR_177 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_9_DFFSR_253 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_36_DFFSR_180 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_26_DFFSR_183 INVX1_67/gnd DFFSR_175/S FILL
XFILL_9_CLKBUF1_10 INVX1_67/gnd DFFSR_201/S FILL
XFILL_48_DFFSR_98 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_8_CLKBUF1_13 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_10_DFFSR_3 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_16_DFFSR_186 BUFX2_99/A DFFSR_92/S FILL
XFILL_6_NAND3X1_105 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_7_CLKBUF1_16 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_32_DFFSR_48 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_21_DFFSR_88 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_4_DFFSR_95 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_4_INVX1_42 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_1_NOR2X1_65 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_6_CLKBUF1_19 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_49_DFFSR_104 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_5_CLKBUF1_22 OR2X2_1/gnd DFFSR_59/S FILL
XNAND3X1_141 NOR2X1_66/Y NAND2X1_64/A NAND2X1_64/B DFFSR_46/gnd AOI21X1_7/B DFFSR_62/S
+ NAND3X1
XFILL_43_1_2 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_39_DFFSR_107 OR2X2_6/gnd DFFSR_92/S FILL
XCLKBUF1_19 BUFX2_3/Y BUFX2_8/gnd DFFSR_1/CLK DFFSR_81/S CLKBUF1
XFILL_4_CLKBUF1_25 INVX1_67/gnd DFFSR_201/S FILL
XFILL_5_9 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_2_DFFSR_183 INVX1_67/gnd DFFSR_175/S FILL
XFILL_3_BUFX2_33 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_29_DFFSR_110 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_43_DFFSR_214 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_3_CLKBUF1_28 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_8_AND2X2_24 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_19_DFFSR_113 BUFX2_99/A DFFSR_92/S FILL
XFILL_33_DFFSR_217 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_2_CLKBUF1_31 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_2_NAND2X1_4 BUFX2_98/A DFFSR_6/S FILL
XFILL_23_DFFSR_220 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_1_CLKBUF1_34 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_4_NAND3X1_201 INVX1_1/gnd DFFSR_53/S FILL
XFILL_40_DFFSR_55 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_1_INVX1_89 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_29_DFFSR_95 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_0_CLKBUF1_37 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_13_DFFSR_223 INVX1_39/gnd DFFSR_34/S FILL
XFILL_0_DFFPOSX1_20 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_11_0_0 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_7_DFFSR_12 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_13_DFFSR_45 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_5_DFFSR_110 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_0_BUFX2_80 BUFX2_79/A DFFSR_6/S FILL
XFILL_2_OAI22X1_3 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_46_DFFSR_141 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_5_NAND3X1_135 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_9_DFFSR_217 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_36_DFFSR_144 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_50_DFFSR_248 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_26_DFFSR_147 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_40_DFFSR_251 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_2_INVX1_194 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_48_DFFSR_62 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_44_5 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_16_DFFSR_150 AND2X2_38/B DFFSR_23/S FILL
XFILL_30_DFFSR_254 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_20_DFFSR_257 INVX1_39/gnd DFFSR_34/S FILL
XFILL_19_DFFPOSX1_28 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_32_DFFSR_12 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_21_DFFSR_52 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_4_DFFSR_59 AND2X2_38/B DFFSR_59/S FILL
XFILL_1_NOR2X1_29 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_10_DFFSR_92 BUFX2_99/A DFFSR_92/S FILL
XFILL_10_DFFSR_260 BUFX2_77/gnd DFFSR_5/S FILL
XNAND3X1_105 DFFSR_190/D BUFX2_29/Y BUFX2_25/Y DFFSR_1/gnd NAND3X1_105/Y DFFSR_81/S
+ NAND3X1
XFILL_3_NAND3X1_231 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_2_DFFSR_147 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_43_DFFSR_178 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_6_DFFSR_254 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_33_DFFSR_181 INVX1_3/gnd DFFSR_79/S FILL
XFILL_23_DFFSR_184 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_4_NAND3X1_165 INVX1_39/gnd DFFSR_34/S FILL
XFILL_40_DFFSR_19 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_1_INVX1_53 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_18_DFFSR_99 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_29_DFFSR_59 AND2X2_38/B DFFSR_59/S FILL
XFILL_13_DFFSR_187 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_9_DFFPOSX1_39 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_0_BUFX2_44 INVX1_3/gnd DFFSR_79/S FILL
XFILL_46_DFFSR_105 INVX1_1/gnd DFFSR_53/S FILL
XFILL_9_DFFSR_181 INVX1_3/gnd DFFSR_79/S FILL
XFILL_36_DFFSR_108 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_50_DFFSR_212 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_26_DFFSR_111 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_40_DFFSR_215 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_2_INVX1_158 INVX1_39/gnd DFFSR_34/S FILL
XFILL_37_DFFSR_66 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_48_DFFSR_26 BUFX2_79/A DFFSR_6/S FILL
XFILL_5_AND2X2_25 INVX1_39/gnd DFFSR_54/S FILL
XFILL_16_DFFSR_114 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_30_DFFSR_218 BUFX2_98/A DFFSR_32/S FILL
XFILL_20_DFFSR_221 AND2X2_38/B DFFSR_59/S FILL
XFILL_21_DFFSR_16 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_4_DFFSR_23 AND2X2_38/B DFFSR_23/S FILL
XFILL_10_DFFSR_56 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_5_OAI21X1_117 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_10_DFFSR_224 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_9_OAI22X1_1 INVX1_1/gnd DFFSR_53/S FILL
XFILL_3_NAND3X1_195 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_2_DFFSR_111 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_3_NOR2X1_4 INVX1_1/gnd DFFSR_53/S FILL
XFILL_43_DFFSR_142 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_22_DFFSR_6 BUFX2_79/A DFFSR_6/S FILL
XFILL_45_DFFSR_73 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_6_DFFSR_218 BUFX2_98/A DFFSR_32/S FILL
XFILL_33_DFFSR_145 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_47_DFFSR_249 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_23_DFFSR_148 INVX1_67/gnd DFFSR_175/S FILL
XFILL_44_2_0 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_4_NAND3X1_129 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_1_DFFSR_70 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_37_DFFSR_252 AND2X2_38/B DFFSR_23/S FILL
XFILL_1_INVX1_17 AND2X2_38/B DFFSR_59/S FILL
XFILL_18_DFFSR_63 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_29_DFFSR_23 AND2X2_38/B DFFSR_23/S FILL
XFILL_13_DFFSR_151 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_5_BUFX2_98 BUFX2_79/A DFFSR_7/S FILL
XFILL_6_BUFX2_7 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_27_DFFSR_255 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_42_4_1 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_6_NAND2X1_165 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_17_DFFSR_258 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_9_DFFSR_145 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_40_6_2 BUFX2_98/A DFFSR_6/S FILL
XFILL_43_DFFSR_2 BUFX2_79/A DFFSR_7/S FILL
XFILL_20_DFFPOSX1_1 INVX1_39/gnd DFFSR_34/S FILL
XFILL_18_DFFPOSX1_22 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_50_DFFSR_176 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_19_DFFPOSX1_4 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_40_DFFSR_179 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_2_INVX1_122 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_26_DFFSR_70 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_37_DFFSR_30 BUFX2_98/A DFFSR_32/S FILL
XFILL_9_DFFSR_77 BUFX2_98/A DFFSR_32/S FILL
XFILL_2_NAND3X1_225 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_18_DFFPOSX1_7 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_3_DFFSR_255 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_30_DFFSR_182 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_20_DFFSR_185 INVX1_39/gnd DFFSR_54/S FILL
XFILL_10_DFFSR_20 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_10_DFFSR_188 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_5_NOR2X1_64 AND2X2_38/B DFFSR_59/S FILL
XFILL_3_NAND3X1_159 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_1_NOR3X1_1 INVX1_3/gnd DFFSR_79/S FILL
XFILL_4_1 INVX1_67/gnd DFFSR_175/S FILL
XFILL_8_DFFPOSX1_33 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_43_DFFSR_106 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_45_DFFSR_37 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_34_DFFSR_77 BUFX2_98/A DFFSR_32/S FILL
XFILL_6_DFFSR_182 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_33_DFFSR_109 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_47_DFFSR_213 INVX1_3/gnd DFFSR_23/S FILL
XFILL_23_DFFSR_112 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_37_DFFSR_216 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_1_DFFSR_34 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_18_DFFSR_27 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_2_AND2X2_26 INVX1_1/gnd DFFSR_97/S FILL
XFILL_6_NAND2X1_3 BUFX2_99/A DFFSR_7/S FILL
XFILL_13_DFFSR_115 INVX1_1/gnd DFFSR_97/S FILL
XFILL_5_BUFX2_62 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_27_DFFSR_219 INVX1_67/gnd DFFSR_175/S FILL
XFILL_10_OAI22X1_8 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_6_NAND2X1_129 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_17_DFFSR_222 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_50_1_2 DFFSR_4/gnd DFFSR_4/S FILL
XXOR2X1_4 XOR2X1_4/A XOR2X1_4/B XOR2X1_4/gnd XOR2X1_4/Y DFFSR_97/S XOR2X1
XFILL_9_DFFSR_109 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_42_DFFSR_84 BUFX2_99/A DFFSR_7/S FILL
XNAND2X1_165 DFFSR_208/S NAND2X1_165/B DFFSR_62/gnd AOI21X1_58/B DFFSR_208/S NAND2X1
XFILL_6_OAI22X1_2 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_4_OAI21X1_111 AND2X2_38/B DFFSR_59/S FILL
XFILL_50_DFFSR_140 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_8_AOI21X1_57 INVX1_67/gnd DFFSR_201/S FILL
XFILL_27_DFFPOSX1_41 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_40_DFFSR_143 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_9_DFFSR_41 BUFX2_98/A DFFSR_6/S FILL
XFILL_7_AOI21X1_60 BUFX2_79/A DFFSR_7/S FILL
XFILL_26_2 AND2X2_38/B DFFSR_23/S FILL
XFILL_26_DFFSR_34 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_2_NAND3X1_189 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_15_DFFSR_74 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_3_DFFSR_219 INVX1_67/gnd DFFSR_175/S FILL
XFILL_30_DFFSR_146 BUFX2_79/A DFFSR_7/S FILL
XFILL_6_AOI21X1_63 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_44_DFFSR_250 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_20_DFFSR_149 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_5_AOI21X1_66 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_34_DFFSR_253 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_18_0_0 DFFSR_1/gnd DFFSR_1/S FILL
XAOI21X1_63 NOR3X1_6/B NOR3X1_6/C AOI21X1_63/C NOR3X1_6/gnd AOI21X1_63/Y DFFSR_91/S
+ AOI21X1
XFILL_10_DFFSR_152 INVX1_1/gnd DFFSR_53/S FILL
XFILL_4_AOI21X1_69 INVX1_1/gnd DFFSR_97/S FILL
XFILL_24_DFFSR_256 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_5_NOR2X1_28 BUFX2_98/A DFFSR_6/S FILL
XFILL_3_NAND3X1_123 BUFX2_99/A DFFSR_7/S FILL
XFILL_50_DFFSR_91 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_14_DFFSR_259 BUFX2_79/A DFFSR_6/S FILL
XFILL_16_2_1 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_5_NAND2X1_159 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_6_DFFSR_88 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_34_DFFSR_41 BUFX2_98/A DFFSR_6/S FILL
XFILL_23_DFFSR_81 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_6_DFFSR_146 BUFX2_79/A DFFSR_7/S FILL
XFILL_14_4_2 INVX1_39/gnd DFFSR_54/S FILL
XFILL_47_DFFSR_177 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_37_DFFSR_180 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_8_OR2X2_5 BUFX2_8/gnd DFFSR_81/S FILL
XBUFX2_66 BUFX2_60/A DFFSR_1/gnd BUFX2_66/Y DFFSR_81/S BUFX2
XFILL_0_DFFSR_256 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_5_BUFX2_26 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_27_DFFSR_183 INVX1_67/gnd DFFSR_175/S FILL
XFILL_17_DFFPOSX1_16 INVX1_67/gnd DFFSR_175/S FILL
XFILL_17_DFFSR_186 BUFX2_99/A DFFSR_92/S FILL
XFILL_15_NOR3X1_5 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_34_DFFSR_9 BUFX2_79/A DFFSR_6/S FILL
XFILL_1_NAND3X1_219 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_3_INVX1_82 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_42_DFFSR_48 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_8_DFFPOSX1_1 INVX1_39/gnd DFFSR_34/S FILL
XFILL_31_DFFSR_88 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_2_NOR2X1_65 DFFSR_34/gnd DFFSR_1/S FILL
XNAND2X1_129 BUFX2_52/Y INVX1_162/A DFFSR_46/gnd OAI21X1_98/C DFFSR_54/S NAND2X1
XFILL_50_DFFSR_104 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_8_AOI21X1_21 INVX1_39/gnd DFFSR_54/S FILL
XFILL_7_DFFPOSX1_4 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_40_DFFSR_107 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_9_6 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_6_DFFPOSX1_7 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_7_AOI21X1_24 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_15_DFFSR_38 BUFX2_98/A DFFSR_6/S FILL
XFILL_2_NAND3X1_153 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_3_DFFSR_183 INVX1_67/gnd DFFSR_175/S FILL
XFILL_30_DFFSR_110 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_2_BUFX2_73 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_6_AOI21X1_27 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_44_DFFSR_214 BUFX2_72/gnd DFFSR_276/S FILL
XDFFPOSX1_7 NOR3X1_4/A CLKBUF1_46/Y OAI21X1_19/Y OR2X2_3/gnd DFFSR_4/S DFFPOSX1
XFILL_20_DFFSR_113 BUFX2_99/A DFFSR_92/S FILL
XFILL_7_DFFPOSX1_27 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_34_DFFSR_217 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_5_AOI21X1_30 XOR2X1_4/gnd DFFSR_97/S FILL
XAOI21X1_27 AOI21X1_27/A AOI21X1_27/B AOI21X1_27/C OR2X2_1/gnd OAI21X1_73/A DFFSR_51/S
+ AOI21X1
XFILL_3_NAND2X1_4 BUFX2_98/A DFFSR_6/S FILL
XFILL_10_DFFSR_116 INVX1_3/gnd DFFSR_23/S FILL
XFILL_4_AOI21X1_33 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_24_DFFSR_220 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_50_DFFSR_55 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_39_DFFSR_95 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_3_AOI21X1_36 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_14_DFFSR_223 INVX1_39/gnd DFFSR_34/S FILL
XFILL_2_AOI21X1_39 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_16_DFFPOSX1_46 INVX1_39/gnd DFFSR_34/S FILL
XFILL_0_AND2X2_4 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_6_DFFSR_52 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_5_NAND2X1_123 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_12_DFFSR_85 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_23_DFFSR_45 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_6_DFFSR_110 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_1_AOI21X1_42 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_3_OAI22X1_3 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_0_NAND3X1_249 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_47_DFFSR_141 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_0_AOI21X1_45 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_37_DFFSR_144 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_51_DFFSR_248 DFFSR_28/gnd DFFSR_8/S FILL
XBUFX2_30 BUFX2_27/A OR2X2_1/gnd BUFX2_30/Y DFFSR_51/S BUFX2
XFILL_4_0_2 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_0_DFFSR_220 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_27_DFFSR_147 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_3_OAI21X1_105 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_41_DFFSR_251 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_26_DFFPOSX1_35 INVX1_39/gnd DFFSR_54/S FILL
XFILL_3_INVX1_194 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_48_2 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_17_DFFSR_150 AND2X2_38/B DFFSR_23/S FILL
XFILL_8_OAI21X1_69 INVX1_3/gnd DFFSR_23/S FILL
XFILL_1_NAND3X1_183 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_31_DFFSR_254 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_7_OAI21X1_72 INVX1_3/gnd DFFSR_23/S FILL
XFILL_6_NAND2X1_90 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_21_DFFSR_257 INVX1_39/gnd DFFSR_34/S FILL
XFILL_42_DFFSR_12 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_31_DFFSR_52 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_3_INVX1_46 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_3_DFFSR_99 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_20_DFFSR_92 BUFX2_99/A DFFSR_92/S FILL
XFILL_2_NOR2X1_29 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_5_NAND2X1_93 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_11_DFFSR_260 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_6_OAI21X1_75 INVX1_39/gnd DFFSR_54/S FILL
XNAND2X1_90 NAND2X1_90/A NAND2X1_90/B DFFSR_46/gnd NAND2X1_90/Y DFFSR_54/S NAND2X1
XFILL_5_OAI21X1_78 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_4_NAND2X1_96 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_51_2_0 DFFSR_4/gnd DFFSR_98/S FILL
XOAI21X1_75 AOI21X1_35/Y OAI21X1_75/B INVX1_131/Y INVX1_39/gnd OAI22X1_51/D DFFSR_54/S
+ OAI21X1
XFILL_2_NAND3X1_117 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_4_OAI21X1_81 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_3_DFFSR_147 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_3_NAND2X1_99 INVX1_39/gnd DFFSR_54/S FILL
XFILL_2_BUFX2_37 INVX1_1/gnd DFFSR_97/S FILL
XFILL_44_DFFSR_178 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_3_OAI21X1_84 BUFX2_98/A DFFSR_6/S FILL
XFILL_7_DFFSR_254 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_49_4_1 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_4_NAND2X1_153 BUFX2_98/A DFFSR_32/S FILL
XFILL_34_DFFSR_181 INVX1_3/gnd DFFSR_79/S FILL
XFILL_21_DFFSR_3 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_2_OAI21X1_87 BUFX2_79/A DFFSR_7/S FILL
XFILL_24_DFFSR_184 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_1_OAI21X1_90 BUFX2_98/A DFFSR_32/S FILL
XFILL_50_DFFSR_19 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_28_DFFSR_99 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_0_INVX1_93 INVX1_3/gnd DFFSR_23/S FILL
XFILL_39_DFFSR_59 AND2X2_38/B DFFSR_59/S FILL
XFILL_47_6_2 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_14_DFFSR_187 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_0_OAI21X1_93 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_16_DFFPOSX1_10 INVX1_67/gnd DFFSR_201/S FILL
XFILL_6_DFFSR_16 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_5_BUFX2_4 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_12_DFFSR_49 OR2X2_6/gnd DFFSR_92/S FILL
XBUFX2_8 BUFX2_7/A BUFX2_8/gnd BUFX2_8/Y DFFSR_51/S BUFX2
XFILL_47_DFFSR_105 INVX1_1/gnd DFFSR_53/S FILL
XFILL_0_NAND3X1_213 INVX1_39/gnd DFFSR_54/S FILL
XFILL_37_DFFSR_108 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_0_DFFSR_184 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_27_DFFSR_111 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_9_OAI21X1_30 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_41_DFFSR_215 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_47_DFFSR_66 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_3_INVX1_158 INVX1_39/gnd DFFSR_34/S FILL
XFILL_6_AND2X2_25 INVX1_39/gnd DFFSR_54/S FILL
XFILL_17_DFFSR_114 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_8_OAI21X1_33 INVX1_3/gnd DFFSR_79/S FILL
XFILL_15_5_0 INVX1_39/gnd DFFSR_34/S FILL
XFILL_31_DFFSR_218 BUFX2_98/A DFFSR_32/S FILL
XFILL_1_NAND3X1_147 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_0_NAND2X1_5 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_6_NAND2X1_54 AND2X2_38/B DFFSR_59/S FILL
XFILL_7_OAI21X1_36 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_21_DFFSR_221 AND2X2_38/B DFFSR_59/S FILL
XFILL_31_DFFSR_16 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_3_DFFSR_63 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_3_INVX1_10 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_20_DFFSR_56 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_6_DFFPOSX1_21 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_5_NAND2X1_57 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_11_DFFSR_224 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_6_OAI21X1_39 DFFSR_34/gnd DFFSR_1/S FILL
XNAND2X1_54 NOR3X1_4/B INVX1_124/Y AND2X2_38/B NAND2X1_54/Y DFFSR_59/S NAND2X1
XFILL_5_OAI21X1_42 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_4_NAND2X1_60 DFFSR_34/gnd DFFSR_34/S FILL
XOAI21X1_39 OAI21X1_41/A OAI21X1_41/B INVX1_152/Y DFFSR_34/gnd AOI22X1_20/C DFFSR_1/S
+ OAI21X1
XFILL_3_DFFSR_111 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_3_NAND2X1_63 AND2X2_38/B DFFSR_59/S FILL
XFILL_4_OAI21X1_45 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_0_OAI22X1_4 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_44_DFFSR_142 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_15_DFFPOSX1_40 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_3_OAI21X1_48 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_2_NAND2X1_66 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_7_DFFSR_218 BUFX2_98/A DFFSR_32/S FILL
XFILL_34_DFFSR_145 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_4_NAND2X1_117 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_48_DFFSR_249 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_1_NAND2X1_69 INVX1_3/gnd DFFSR_23/S FILL
XFILL_2_OAI21X1_51 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_24_DFFSR_148 INVX1_67/gnd DFFSR_175/S FILL
XFILL_38_DFFSR_252 AND2X2_38/B DFFSR_23/S FILL
XFILL_0_NAND2X1_72 AND2X2_38/B DFFSR_59/S FILL
XFILL_1_OAI21X1_54 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_28_DFFSR_63 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_0_INVX1_57 BUFX2_98/A DFFSR_32/S FILL
XFILL_39_DFFSR_23 AND2X2_38/B DFFSR_23/S FILL
XFILL_10_AOI22X1_20 INVX1_39/gnd DFFSR_34/S FILL
XFILL_0_INVX1_195 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_14_DFFSR_151 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_0_OAI21X1_57 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_28_DFFSR_255 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_25_DFFPOSX1_29 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_18_DFFSR_258 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_12_DFFSR_13 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_9_AOI22X1_23 INVX1_39/gnd DFFSR_34/S FILL
XFILL_8_AOI22X1_26 INVX1_1/gnd DFFSR_97/S FILL
XFILL_0_NAND3X1_177 AND2X2_38/B DFFSR_59/S FILL
XFILL_9_NAND3X1_232 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_7_AOI22X1_29 INVX1_1/gnd DFFSR_53/S FILL
XNOR2X1_1 BUFX2_8/Y INVX1_4/Y BUFX2_99/A NOR2X1_1/Y DFFSR_92/S NOR2X1
XFILL_51_DFFSR_176 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_0_DFFSR_148 INVX1_67/gnd DFFSR_175/S FILL
XDFFSR_258 DFFSR_2/D CLKBUF1_4/Y DFFSR_257/R DFFSR_5/S DFFSR_258/D DFFSR_5/gnd DFFSR_5/S
+ DFFSR
XFILL_25_0_0 AND2X2_38/B DFFSR_23/S FILL
XFILL_41_DFFSR_179 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_47_DFFSR_30 BUFX2_98/A DFFSR_32/S FILL
XFILL_3_INVX1_122 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_36_DFFSR_70 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_4_DFFSR_255 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_31_DFFSR_182 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_1_NAND3X1_111 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_23_2_1 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_6_NAND2X1_18 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_21_DFFSR_185 INVX1_39/gnd DFFSR_54/S FILL
XFILL_3_DFFSR_27 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_20_DFFSR_20 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_5_1_0 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_5_NAND2X1_21 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_3_NAND2X1_147 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_11_DFFSR_188 DFFSR_46/gnd DFFSR_54/S FILL
XNAND2X1_18 DFFSR_44/D AND2X2_5/Y OR2X2_3/gnd NAND3X1_28/A DFFSR_60/S NAND2X1
XFILL_21_4_2 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_4_NAND2X1_24 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_6_NOR2X1_64 AND2X2_38/B DFFSR_59/S FILL
XFILL_3_3_1 INVX1_67/gnd DFFSR_175/S FILL
XFILL_9_DFFSR_2 BUFX2_79/A DFFSR_7/S FILL
XFILL_2_NOR2X1_8 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_3_NAND2X1_27 AND2X2_38/B DFFSR_23/S FILL
XDFFPOSX1_21 INVX1_180/A CLKBUF1_46/Y NAND2X1_115/Y DFFSR_28/gnd DFFSR_8/S DFFPOSX1
XFILL_44_DFFSR_106 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_2_NAND2X1_30 AND2X2_38/B DFFSR_23/S FILL
XFILL_3_OAI21X1_12 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_44_DFFSR_77 BUFX2_98/A DFFSR_32/S FILL
XFILL_7_DFFSR_182 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_34_DFFSR_109 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_1_NAND2X1_33 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_2_OAI21X1_15 INVX1_3/gnd DFFSR_79/S FILL
XFILL_48_DFFSR_213 INVX1_3/gnd DFFSR_23/S FILL
XFILL_1_5_2 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_24_DFFSR_112 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_8_NAND3X1_89 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_38_DFFSR_216 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_0_NAND2X1_36 INVX1_3/gnd DFFSR_79/S FILL
XFILL_1_OAI21X1_18 INVX1_39/gnd DFFSR_34/S FILL
XFILL_28_DFFSR_27 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_0_DFFSR_74 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_0_INVX1_21 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_0_INVX1_159 INVX1_3/gnd DFFSR_79/S FILL
XFILL_17_DFFSR_67 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_3_AND2X2_26 INVX1_1/gnd DFFSR_97/S FILL
XFILL_14_DFFSR_115 INVX1_1/gnd DFFSR_97/S FILL
XFILL_7_NAND3X1_92 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_0_OAI21X1_21 AND2X2_38/B DFFSR_59/S FILL
XFILL_28_DFFSR_219 INVX1_67/gnd DFFSR_175/S FILL
XFILL_11_OAI22X1_8 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_6_NAND3X1_95 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_7_OR2X2_2 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_18_DFFSR_222 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_5_NAND3X1_98 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_4_XOR2X1_4 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_0_NAND3X1_141 DFFSR_46/gnd DFFSR_62/S FILL
XNAND3X1_95 NAND3X1_93/Y NAND3X1_94/Y AOI22X1_12/Y DFFSR_62/gnd NOR2X1_46/B DFFSR_208/S
+ NAND3X1
XFILL_33_DFFSR_6 BUFX2_79/A DFFSR_6/S FILL
XFILL_7_OAI22X1_2 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_5_DFFPOSX1_15 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_51_DFFSR_140 DFFSR_62/gnd DFFSR_208/S FILL
XDFFSR_222 DFFSR_222/Q CLKBUF1_25/Y BUFX2_60/Y DFFSR_201/S INVX1_99/A BUFX2_72/gnd
+ DFFSR_201/S DFFSR
XFILL_0_DFFSR_112 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_2_NAND2X1_177 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_41_DFFSR_143 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_8_DFFSR_81 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_36_DFFSR_34 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_25_DFFSR_74 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_4_DFFSR_219 INVX1_67/gnd DFFSR_175/S FILL
XFILL_31_DFFSR_146 BUFX2_79/A DFFSR_7/S FILL
XFILL_45_DFFSR_250 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_21_DFFSR_149 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_14_DFFPOSX1_34 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_35_DFFSR_253 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_3_NAND2X1_111 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_11_DFFSR_152 INVX1_1/gnd DFFSR_53/S FILL
XFILL_25_DFFSR_256 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_6_NOR2X1_28 BUFX2_98/A DFFSR_6/S FILL
XFILL_15_DFFSR_259 BUFX2_79/A DFFSR_6/S FILL
XFILL_0_NOR3X1_5 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_1_AOI22X1_11 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_0_AOI22X1_14 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_10_OAI22X1_32 INVX1_39/gnd DFFSR_54/S FILL
XFILL_44_DFFSR_41 BUFX2_98/A DFFSR_6/S FILL
XFILL_33_DFFSR_81 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_7_DFFSR_146 BUFX2_79/A DFFSR_7/S FILL
XFILL_24_DFFPOSX1_23 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_48_DFFSR_177 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_8_NAND3X1_53 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_9_OAI22X1_35 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_38_DFFSR_180 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_8_NAND3X1_226 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_0_DFFSR_38 BUFX2_98/A DFFSR_6/S FILL
XFILL_17_DFFSR_31 BUFX2_79/A DFFSR_6/S FILL
XFILL_0_INVX1_123 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_7_NAND3X1_56 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_1_DFFSR_256 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_8_OAI22X1_38 AND2X2_38/B DFFSR_23/S FILL
XFILL_4_BUFX2_66 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_28_DFFSR_183 INVX1_67/gnd DFFSR_175/S FILL
XFILL_4_DFFPOSX1_45 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_6_NAND3X1_59 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_7_OAI22X1_41 INVX1_39/gnd DFFSR_54/S FILL
XFILL_18_DFFSR_186 BUFX2_99/A DFFSR_92/S FILL
XFILL_5_NAND3X1_62 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_6_OAI22X1_44 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_0_NAND3X1_105 DFFSR_1/gnd DFFSR_81/S FILL
XNAND3X1_59 BUFX2_89/A AND2X2_3/Y BUFX2_21/Y OR2X2_4/gnd AND2X2_13/A DFFSR_32/S NAND3X1
XFILL_10_XOR2X1_1 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_5_OAI22X1_47 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_4_NAND3X1_65 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_41_DFFSR_88 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_3_NOR2X1_65 DFFSR_34/gnd DFFSR_1/S FILL
XOAI22X1_44 INVX1_106/Y OAI22X1_41/B INVX1_107/Y OAI22X1_41/D DFFSR_1/gnd NOR2X1_53/A
+ DFFSR_81/S OAI22X1
XFILL_3_NAND3X1_68 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_4_OAI22X1_50 INVX1_3/gnd DFFSR_23/S FILL
XDFFSR_186 INVX1_70/A CLKBUF1_3/Y BUFX2_63/Y DFFSR_92/S DFFSR_170/Q BUFX2_99/A DFFSR_92/S
+ DFFSR
XFILL_2_NAND2X1_141 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_2_NAND3X1_71 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_41_DFFSR_107 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_8_DFFSR_45 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_14_DFFSR_78 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_25_DFFSR_38 BUFX2_98/A DFFSR_6/S FILL
XFILL_4_DFFSR_183 INVX1_67/gnd DFFSR_175/S FILL
XFILL_31_DFFSR_110 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_1_NAND3X1_74 INVX1_1/gnd DFFSR_97/S FILL
XFILL_45_DFFSR_214 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_54_6_2 DFFSR_5/gnd DFFSR_5/S FILL
XNAND2X1_7 BUFX2_9/Y INVX1_4/Y OR2X2_6/gnd NOR2X1_5/B DFFSR_53/S NAND2X1
XFILL_0_NAND3X1_77 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_21_DFFSR_113 BUFX2_99/A DFFSR_92/S FILL
XFILL_35_DFFSR_217 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_0_AND2X2_27 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_11_DFFSR_116 INVX1_3/gnd DFFSR_23/S FILL
XFILL_4_NAND2X1_4 BUFX2_98/A DFFSR_6/S FILL
XFILL_25_DFFSR_220 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_0_DFFSR_9 BUFX2_79/A DFFSR_6/S FILL
XFILL_49_DFFSR_95 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_15_DFFSR_223 INVX1_39/gnd DFFSR_34/S FILL
XOAI22X1_6 INVX1_14/Y OAI22X1_6/B INVX1_15/Y OAI22X1_6/D BUFX2_98/A OAI22X1_6/Y DFFSR_32/S
+ OAI22X1
XINVX1_79 INVX1_79/A INVX1_39/gnd INVX1_79/Y DFFSR_54/S INVX1
XFILL_33_DFFSR_45 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_5_DFFSR_92 BUFX2_99/A DFFSR_92/S FILL
XFILL_22_DFFSR_85 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_7_DFFSR_110 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_4_OAI22X1_3 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_48_DFFSR_141 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_22_5_0 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_4_BUFX2_1 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_8_NAND3X1_17 BUFX2_99/A DFFSR_7/S FILL
XFILL_38_DFFSR_144 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_8_NAND3X1_190 BUFX2_7/gnd DFFSR_151/S FILL
XINVX1_197 DFFSR_272/Q INVX1_3/gnd INVX1_197/Y DFFSR_79/S INVX1
XFILL_1_DFFSR_220 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_7_NAND3X1_20 BUFX2_99/A DFFSR_7/S FILL
XFILL_4_BUFX2_30 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_28_DFFSR_147 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_42_DFFSR_251 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_1_NAND2X1_171 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_6_NAND3X1_23 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_18_DFFSR_150 AND2X2_38/B DFFSR_23/S FILL
XFILL_32_DFFSR_254 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_2_6_0 INVX1_67/gnd DFFSR_201/S FILL
XFILL_5_NAND3X1_26 DFFSR_28/gnd DFFSR_3/S FILL
XNAND3X1_23 NAND3X1_23/A NAND3X1_22/Y AOI22X1_3/Y OR2X2_6/gnd NOR2X1_14/B DFFSR_53/S
+ NAND3X1
XFILL_22_DFFSR_257 INVX1_39/gnd DFFSR_34/S FILL
XFILL_4_NAND3X1_29 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_5_OAI22X1_11 BUFX2_99/A DFFSR_92/S FILL
XFILL_41_DFFSR_52 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_30_DFFSR_92 BUFX2_99/A DFFSR_92/S FILL
XFILL_2_INVX1_86 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_3_NOR2X1_29 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_13_DFFPOSX1_28 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_12_DFFSR_260 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_4_OAI22X1_14 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_3_NAND3X1_32 BUFX2_79/A DFFSR_7/S FILL
XFILL_2_NAND2X1_105 OR2X2_6/gnd DFFSR_53/S FILL
XDFFSR_150 INVX1_101/A CLKBUF1_22/Y BUFX2_61/Y DFFSR_23/S INVX1_102/A AND2X2_38/B
+ DFFSR_23/S DFFSR
XFILL_2_NAND3X1_35 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_3_OAI22X1_17 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_14_DFFSR_42 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_4_DFFSR_147 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_1_BUFX2_77 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_2_OAI22X1_20 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_1_NAND3X1_38 BUFX2_98/A DFFSR_32/S FILL
XFILL_45_DFFSR_178 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_1_OAI22X1_23 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_0_NAND3X1_41 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_8_DFFSR_254 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_35_DFFSR_181 INVX1_3/gnd DFFSR_79/S FILL
XFILL_23_DFFPOSX1_17 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_0_OAI22X1_26 INVX1_39/gnd DFFSR_54/S FILL
XFILL_45_DFFSR_9 BUFX2_79/A DFFSR_6/S FILL
XFILL_25_DFFSR_184 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_38_DFFSR_99 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_49_DFFSR_59 AND2X2_38/B DFFSR_59/S FILL
XFILL_15_DFFSR_187 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_7_NAND3X1_220 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_3_DFFPOSX1_39 BUFX2_7/gnd DFFSR_151/S FILL
XINVX1_43 DFFSR_30/Q OR2X2_4/gnd INVX1_43/Y DFFSR_3/S INVX1
XDFFSR_96 DFFSR_96/Q DFFSR_85/CLK DFFSR_5/R DFFSR_4/S INVX1_54/A DFFSR_4/gnd DFFSR_4/S
+ DFFSR
XFILL_32_0_0 INVX1_1/gnd DFFSR_97/S FILL
XFILL_5_DFFSR_56 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_22_DFFSR_49 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_11_DFFSR_89 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_0_NOR2X1_66 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_48_DFFSR_105 INVX1_1/gnd DFFSR_53/S FILL
XFILL_38_DFFSR_108 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_30_2_1 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_8_NAND3X1_154 BUFX2_7/gnd DFFSR_216/S FILL
XINVX1_161 AND2X2_37/B INVX1_1/gnd INVX1_161/Y DFFSR_53/S INVX1
XFILL_1_DFFSR_184 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_28_DFFSR_111 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_42_DFFSR_215 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_1_NAND2X1_135 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_4_INVX1_158 INVX1_39/gnd DFFSR_34/S FILL
XFILL_7_AND2X2_25 INVX1_39/gnd DFFSR_54/S FILL
XFILL_18_DFFSR_114 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_28_4_2 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_32_DFFSR_218 BUFX2_98/A DFFSR_32/S FILL
XFILL_1_NAND2X1_5 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_22_DFFSR_221 AND2X2_38/B DFFSR_59/S FILL
XFILL_2_INVX1_50 BUFX2_98/A DFFSR_6/S FILL
XFILL_41_DFFSR_16 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_30_DFFSR_56 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_19_DFFSR_96 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_12_DFFSR_224 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_22_DFFPOSX1_47 XOR2X1_4/gnd DFFSR_91/S FILL
XDFFSR_114 INVX1_16/A CLKBUF1_27/Y BUFX2_49/Y DFFSR_91/S DFFSR_114/D NOR3X1_6/gnd
+ DFFSR_91/S DFFSR
XFILL_8_5_2 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_4_DFFSR_111 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_1_BUFX2_41 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_1_OAI22X1_4 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_45_DFFSR_142 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_8_DFFSR_218 BUFX2_98/A DFFSR_32/S FILL
XFILL_35_DFFSR_145 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_49_DFFSR_249 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_11_DFFSR_7 BUFX2_79/A DFFSR_7/S FILL
XFILL_25_DFFSR_148 INVX1_67/gnd DFFSR_175/S FILL
XFILL_38_DFFSR_63 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_49_DFFSR_23 AND2X2_38/B DFFSR_23/S FILL
XFILL_39_DFFSR_252 AND2X2_38/B DFFSR_23/S FILL
XFILL_1_INVX1_195 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_15_DFFSR_151 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_7_NAND3X1_184 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_29_DFFSR_255 OR2X2_4/gnd DFFSR_32/S FILL
XDFFSR_60 INVX1_25/A CLKBUF1_4/Y DFFSR_8/R DFFSR_60/S DFFSR_60/D OR2X2_3/gnd DFFSR_60/S
+ DFFSR
XFILL_19_DFFSR_258 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_0_NAND2X1_165 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_5_DFFSR_20 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_22_DFFSR_13 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_11_DFFSR_53 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_0_NOR2X1_30 INVX1_3/gnd DFFSR_23/S FILL
XFILL_8_NAND3X1_118 DFFSR_62/gnd DFFSR_62/S FILL
XINVX1_125 NOR3X1_4/B AND2X2_38/B INVX1_125/Y DFFSR_59/S INVX1
XFILL_1_DFFSR_148 INVX1_67/gnd DFFSR_175/S FILL
XFILL_4_NOR2X1_1 BUFX2_99/A DFFSR_92/S FILL
XFILL_12_DFFPOSX1_22 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_32_DFFSR_3 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_42_DFFSR_179 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_4_INVX1_122 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_46_DFFSR_70 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_5_DFFSR_255 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_32_DFFSR_182 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_22_DFFSR_185 INVX1_39/gnd DFFSR_54/S FILL
XFILL_2_INVX1_14 BUFX2_98/A DFFSR_6/S FILL
XFILL_19_DFFSR_60 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_30_DFFSR_20 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_2_DFFSR_67 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_6_BUFX2_95 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_12_DFFSR_188 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_22_DFFPOSX1_11 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_6_NAND3X1_214 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_45_DFFSR_106 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_2_DFFPOSX1_33 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_8_DFFSR_182 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_35_DFFSR_109 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_49_DFFSR_213 INVX1_3/gnd DFFSR_23/S FILL
XAND2X2_29 BUFX2_59/Y INVX1_145/A AND2X2_38/B AND2X2_29/Y DFFSR_23/S AND2X2
XFILL_25_DFFSR_112 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_39_DFFSR_216 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_38_DFFSR_27 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_1_INVX1_159 INVX1_3/gnd DFFSR_79/S FILL
XFILL_4_AND2X2_26 INVX1_1/gnd DFFSR_97/S FILL
XFILL_27_DFFSR_67 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_15_DFFSR_115 INVX1_1/gnd DFFSR_97/S FILL
XFILL_7_NAND3X1_148 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_29_DFFSR_219 INVX1_67/gnd DFFSR_175/S FILL
XFILL_19_DFFSR_222 BUFX2_72/gnd DFFSR_201/S FILL
XDFFSR_24 DFFSR_24/Q DFFSR_2/CLK DFFSR_2/R DFFSR_6/S DFFSR_24/D BUFX2_98/A DFFSR_6/S
+ DFFSR
XFILL_0_NAND2X1_129 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_11_DFFSR_17 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_8_OAI22X1_2 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_1_DFFSR_112 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_17_1 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_42_DFFSR_143 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_21_DFFPOSX1_41 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_35_DFFSR_74 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_46_DFFSR_34 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_5_DFFSR_219 INVX1_67/gnd DFFSR_175/S FILL
XFILL_32_DFFSR_146 BUFX2_79/A DFFSR_7/S FILL
XFILL_46_DFFSR_250 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_5_NAND3X1_244 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_22_DFFSR_149 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_19_DFFSR_24 BUFX2_98/A DFFSR_6/S FILL
XFILL_2_DFFSR_31 BUFX2_79/A DFFSR_6/S FILL
XFILL_36_DFFSR_253 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_12_DFFSR_152 INVX1_1/gnd DFFSR_53/S FILL
XFILL_6_BUFX2_59 AND2X2_38/B DFFSR_23/S FILL
XFILL_26_DFFSR_256 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_8_OAI21X1_100 INVX1_3/gnd DFFSR_79/S FILL
XFILL_29_5_0 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_16_DFFSR_259 BUFX2_79/A DFFSR_6/S FILL
XFILL_6_NAND3X1_178 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_20_CLKBUF1_14 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_19_CLKBUF1_17 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_43_DFFSR_81 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_8_DFFSR_146 BUFX2_79/A DFFSR_7/S FILL
XFILL_18_CLKBUF1_20 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_49_DFFSR_177 DFFSR_46/gnd DFFSR_54/S FILL
XNAND3X1_214 NAND3X1_214/A NAND3X1_214/B AOI21X1_33/Y DFFSR_46/gnd NAND3X1_219/B DFFSR_62/S
+ NAND3X1
XFILL_9_6_0 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_39_DFFSR_180 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_17_CLKBUF1_23 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_1_INVX1_123 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_27_DFFSR_31 BUFX2_79/A DFFSR_6/S FILL
XFILL_16_DFFSR_71 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_2_DFFSR_256 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_7_NAND3X1_112 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_29_DFFSR_183 INVX1_67/gnd DFFSR_175/S FILL
XFILL_16_CLKBUF1_26 INVX1_1/gnd DFFSR_53/S FILL
XFILL_11_DFFPOSX1_16 INVX1_67/gnd DFFSR_175/S FILL
XFILL_19_DFFSR_186 BUFX2_99/A DFFSR_92/S FILL
XFILL_15_CLKBUF1_29 XOR2X1_4/gnd DFFSR_91/S FILL
XNOR2X1_68 AND2X2_30/B NOR2X1_67/Y OR2X2_2/gnd NOR2X1_68/Y DFFSR_175/S NOR2X1
XFILL_14_CLKBUF1_32 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_3_XOR2X1_8 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_13_CLKBUF1_35 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_4_NOR2X1_65 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_12_CLKBUF1_38 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_42_DFFSR_107 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_11_CLKBUF1_41 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_7_DFFSR_85 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_24_DFFSR_78 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_35_DFFSR_38 BUFX2_98/A DFFSR_6/S FILL
XFILL_5_DFFSR_183 INVX1_67/gnd DFFSR_175/S FILL
XFILL_32_DFFSR_110 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_46_DFFSR_214 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_10_CLKBUF1_44 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_5_NAND3X1_208 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_22_DFFSR_113 BUFX2_99/A DFFSR_92/S FILL
XFILL_36_DFFSR_217 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_1_DFFPOSX1_27 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_39_0_0 BUFX2_79/A DFFSR_6/S FILL
XFILL_1_AND2X2_27 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_6_BUFX2_23 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_12_DFFSR_116 INVX1_3/gnd DFFSR_23/S FILL
XFILL_5_NAND2X1_4 BUFX2_98/A DFFSR_6/S FILL
XFILL_26_DFFSR_220 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_9_CLKBUF1_47 BUFX2_98/A DFFSR_32/S FILL
XFILL_16_DFFSR_223 INVX1_39/gnd DFFSR_34/S FILL
XFILL_44_DFFSR_6 BUFX2_79/A DFFSR_6/S FILL
XFILL_37_2_1 BUFX2_99/A DFFSR_7/S FILL
XFILL_16_NOR3X1_2 INVX1_1/gnd DFFSR_53/S FILL
XFILL_6_NAND3X1_142 INVX1_67/gnd DFFSR_175/S FILL
XFILL_10_DFFPOSX1_46 INVX1_39/gnd DFFSR_34/S FILL
XFILL_43_DFFSR_45 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_32_DFFSR_85 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_8_DFFSR_110 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_5_OAI22X1_3 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_35_4_2 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_49_DFFSR_141 XOR2X1_4/gnd DFFSR_91/S FILL
XNAND3X1_178 INVX1_160/A AOI21X1_30/B NAND2X1_85/Y NOR3X1_6/gnd AOI21X1_27/A DFFSR_91/S
+ NAND3X1
XFILL_39_DFFSR_144 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_16_DFFSR_35 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_22_6 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_2_DFFSR_220 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_3_BUFX2_70 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_39_1 BUFX2_79/A DFFSR_7/S FILL
XFILL_29_DFFSR_147 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_43_DFFSR_251 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_20_DFFPOSX1_35 INVX1_39/gnd DFFSR_54/S FILL
XFILL_19_DFFSR_150 AND2X2_38/B DFFSR_23/S FILL
XFILL_33_DFFSR_254 DFFSR_34/gnd DFFSR_1/S FILL
XNOR2X1_32 NOR2X1_32/A NOR2X1_32/B DFFSR_34/gnd NOR2X1_32/Y DFFSR_34/S NOR2X1
XFILL_4_NAND3X1_238 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_23_DFFSR_257 INVX1_39/gnd DFFSR_34/S FILL
XFILL_40_DFFSR_92 BUFX2_99/A DFFSR_92/S FILL
XFILL_4_NOR2X1_29 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_13_DFFSR_260 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_1_AND2X2_1 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_24_DFFSR_42 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_7_DFFSR_49 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_13_DFFSR_82 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_5_DFFSR_147 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_46_DFFSR_178 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_5_NAND3X1_172 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_9_DFFSR_254 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_36_DFFSR_181 INVX1_3/gnd DFFSR_79/S FILL
XFILL_26_DFFSR_184 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_9_CLKBUF1_11 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_48_DFFSR_99 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_10_DFFSR_4 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_16_DFFSR_187 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_8_CLKBUF1_14 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_6_NAND3X1_106 INVX1_3/gnd DFFSR_23/S FILL
XFILL_7_CLKBUF1_17 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_10_DFFPOSX1_10 INVX1_67/gnd DFFSR_201/S FILL
XFILL_4_DFFSR_96 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_32_DFFSR_49 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_21_DFFSR_89 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_6_CLKBUF1_20 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_1_NOR2X1_66 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_49_DFFSR_105 INVX1_1/gnd DFFSR_53/S FILL
XFILL_5_CLKBUF1_23 DFFSR_4/gnd DFFSR_98/S FILL
XNAND3X1_142 AOI21X1_7/C AOI21X1_7/B AOI21X1_7/A INVX1_67/gnd INVX1_141/A DFFSR_175/S
+ NAND3X1
XFILL_39_DFFSR_108 OR2X2_6/gnd DFFSR_92/S FILL
XCLKBUF1_20 BUFX2_5/Y BUFX2_8/gnd CLKBUF1_20/Y DFFSR_51/S CLKBUF1
XFILL_4_CLKBUF1_26 INVX1_1/gnd DFFSR_53/S FILL
XFILL_2_DFFSR_184 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_3_BUFX2_34 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_29_DFFSR_111 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_3_CLKBUF1_29 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_43_DFFSR_215 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_8_AND2X2_25 INVX1_39/gnd DFFSR_54/S FILL
XFILL_19_DFFSR_114 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_33_DFFSR_218 BUFX2_98/A DFFSR_32/S FILL
XFILL_2_CLKBUF1_32 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_2_NAND2X1_5 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_4_NAND3X1_202 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_23_DFFSR_221 AND2X2_38/B DFFSR_59/S FILL
XFILL_1_CLKBUF1_35 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_40_DFFSR_56 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_29_DFFSR_96 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_1_INVX1_90 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_13_DFFSR_224 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_0_DFFPOSX1_21 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_0_CLKBUF1_38 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_11_0_1 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_7_DFFSR_13 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_13_DFFSR_46 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_5_DFFSR_111 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_2_OAI22X1_4 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_0_BUFX2_81 BUFX2_79/A DFFSR_7/S FILL
XFILL_46_DFFSR_142 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_5_NAND3X1_136 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_9_DFFSR_218 BUFX2_98/A DFFSR_32/S FILL
XFILL_36_DFFSR_145 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_50_DFFSR_249 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_26_DFFSR_148 INVX1_67/gnd DFFSR_175/S FILL
XFILL_48_DFFSR_63 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_40_DFFSR_252 AND2X2_38/B DFFSR_23/S FILL
XFILL_2_INVX1_195 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_16_DFFSR_151 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_44_6 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_30_DFFSR_255 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_20_DFFSR_258 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_4_DFFSR_60 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_19_DFFPOSX1_29 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_10_DFFSR_93 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_32_DFFSR_13 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_21_DFFSR_53 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_1_NOR2X1_30 INVX1_3/gnd DFFSR_23/S FILL
XFILL_10_DFFSR_261 BUFX2_77/gnd DFFSR_98/S FILL
XNAND3X1_106 DFFSR_158/D AND2X2_18/B BUFX2_29/Y INVX1_3/gnd AND2X2_24/B DFFSR_23/S
+ NAND3X1
XFILL_3_NAND3X1_232 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_2_DFFSR_148 INVX1_67/gnd DFFSR_175/S FILL
XFILL_43_DFFSR_179 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_6_DFFSR_255 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_36_5_0 BUFX2_99/A DFFSR_92/S FILL
XFILL_33_DFFSR_182 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_4_NAND3X1_166 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_23_DFFSR_185 INVX1_39/gnd DFFSR_54/S FILL
XFILL_29_DFFSR_60 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_1_INVX1_54 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_40_DFFSR_20 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_13_DFFSR_188 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_9_DFFPOSX1_40 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_13_DFFSR_10 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_0_BUFX2_45 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_46_DFFSR_106 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_5_NAND3X1_100 AND2X2_38/B DFFSR_59/S FILL
XFILL_9_DFFSR_182 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_36_DFFSR_109 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_50_DFFSR_213 INVX1_3/gnd DFFSR_23/S FILL
XFILL_26_DFFSR_112 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_40_DFFSR_216 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_48_DFFSR_27 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_2_INVX1_159 INVX1_3/gnd DFFSR_79/S FILL
XFILL_5_AND2X2_26 INVX1_1/gnd DFFSR_97/S FILL
XFILL_37_DFFSR_67 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_16_DFFSR_115 INVX1_1/gnd DFFSR_97/S FILL
XFILL_30_DFFSR_219 INVX1_67/gnd DFFSR_175/S FILL
XFILL_20_DFFSR_222 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_4_DFFSR_24 BUFX2_98/A DFFSR_6/S FILL
XFILL_21_DFFSR_17 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_10_DFFSR_57 BUFX2_79/A DFFSR_6/S FILL
XFILL_5_OAI21X1_118 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_10_DFFSR_225 INVX1_67/gnd DFFSR_175/S FILL
XFILL_3_NAND3X1_196 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_9_OAI22X1_2 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_2_DFFSR_112 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_3_NOR2X1_5 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_46_0_0 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_43_DFFSR_143 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_22_DFFSR_7 BUFX2_79/A DFFSR_7/S FILL
XFILL_45_DFFSR_74 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_6_DFFSR_219 INVX1_67/gnd DFFSR_175/S FILL
XFILL_33_DFFSR_146 BUFX2_79/A DFFSR_7/S FILL
XFILL_47_DFFSR_250 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_44_2_1 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_23_DFFSR_149 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_4_NAND3X1_130 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_29_DFFSR_24 BUFX2_98/A DFFSR_6/S FILL
XFILL_1_DFFSR_71 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_1_INVX1_18 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_37_DFFSR_253 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_18_DFFSR_64 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_13_DFFSR_152 INVX1_1/gnd DFFSR_53/S FILL
XFILL_5_BUFX2_99 BUFX2_99/A DFFSR_7/S FILL
XFILL_27_DFFSR_256 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_6_BUFX2_8 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_42_4_2 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_6_NAND2X1_166 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_17_DFFSR_259 BUFX2_79/A DFFSR_6/S FILL
XFILL_5_XOR2X1_1 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_43_DFFSR_3 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_9_DFFSR_146 BUFX2_79/A DFFSR_7/S FILL
XFILL_20_DFFPOSX1_2 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_18_DFFPOSX1_23 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_50_DFFSR_177 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_19_DFFPOSX1_5 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_9_DFFSR_78 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_2_INVX1_123 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_40_DFFSR_180 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_37_DFFSR_31 BUFX2_79/A DFFSR_6/S FILL
XFILL_26_DFFSR_71 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_3_DFFSR_256 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_2_NAND3X1_226 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_18_DFFPOSX1_8 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_30_DFFSR_183 INVX1_67/gnd DFFSR_175/S FILL
XFILL_10_3_0 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_20_DFFSR_186 BUFX2_99/A DFFSR_92/S FILL
XFILL_10_DFFSR_21 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_10_DFFSR_189 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_3_NAND3X1_160 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_5_NOR2X1_65 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_1_NOR3X1_2 INVX1_1/gnd DFFSR_53/S FILL
XFILL_43_DFFSR_107 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_8_DFFPOSX1_34 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_34_DFFSR_78 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_45_DFFSR_38 BUFX2_98/A DFFSR_6/S FILL
XFILL_6_DFFSR_183 INVX1_67/gnd DFFSR_175/S FILL
XFILL_33_DFFSR_110 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_47_DFFSR_214 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_23_DFFSR_113 BUFX2_99/A DFFSR_92/S FILL
XFILL_37_DFFSR_217 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_1_DFFSR_35 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_18_DFFSR_28 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_2_AND2X2_27 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_13_DFFSR_116 INVX1_3/gnd DFFSR_23/S FILL
XFILL_5_BUFX2_63 BUFX2_98/A DFFSR_32/S FILL
XFILL_6_NAND2X1_4 BUFX2_98/A DFFSR_6/S FILL
XFILL_27_DFFSR_220 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_10_OAI22X1_9 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_6_NAND2X1_130 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_17_DFFSR_223 INVX1_39/gnd DFFSR_34/S FILL
XXOR2X1_5 XOR2X1_5/A XOR2X1_5/B OR2X2_6/gnd XOR2X1_5/Y DFFSR_92/S XOR2X1
XFILL_42_DFFSR_85 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_9_DFFSR_110 OR2X2_3/gnd DFFSR_4/S FILL
XNAND2X1_166 NAND2X1_165/B INVX1_208/Y BUFX2_8/gnd AOI21X1_59/A DFFSR_81/S NAND2X1
XFILL_6_OAI22X1_3 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_50_DFFSR_141 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_8_AOI21X1_58 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_4_OAI21X1_112 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_27_DFFPOSX1_42 INVX1_39/gnd DFFSR_34/S FILL
XFILL_9_DFFSR_42 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_40_DFFSR_144 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_26_DFFSR_35 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_7_AOI21X1_61 AND2X2_38/B DFFSR_59/S FILL
XFILL_15_DFFSR_75 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_3_DFFSR_220 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_2_NAND3X1_190 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_30_DFFSR_147 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_6_AOI21X1_64 AND2X2_38/B DFFSR_59/S FILL
XFILL_44_DFFSR_251 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_20_DFFSR_150 AND2X2_38/B DFFSR_23/S FILL
XFILL_5_AOI21X1_67 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_18_0_1 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_34_DFFSR_254 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_10_DFFSR_153 INVX1_67/gnd DFFSR_201/S FILL
XAOI21X1_64 AOI21X1_64/A XOR2X1_10/Y AOI21X1_64/C AND2X2_38/B AOI21X1_64/Y DFFSR_59/S
+ AOI21X1
XFILL_4_AOI21X1_70 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_24_DFFSR_257 INVX1_39/gnd DFFSR_34/S FILL
XFILL_50_DFFSR_92 BUFX2_99/A DFFSR_92/S FILL
XFILL_5_NOR2X1_29 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_3_NAND3X1_124 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_14_DFFSR_260 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_16_2_2 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_34_DFFSR_42 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_5_NAND2X1_160 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_6_DFFSR_89 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_23_DFFSR_82 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_6_DFFSR_147 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_47_DFFSR_178 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_37_DFFSR_181 INVX1_3/gnd DFFSR_79/S FILL
XFILL_8_OR2X2_6 OR2X2_6/gnd DFFSR_53/S FILL
XBUFX2_67 BUFX2_60/A OR2X2_2/gnd BUFX2_67/Y DFFSR_216/S BUFX2
XFILL_0_DFFSR_257 INVX1_39/gnd DFFSR_34/S FILL
XFILL_5_BUFX2_27 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_27_DFFSR_184 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_17_DFFPOSX1_17 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_17_DFFSR_187 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_15_NOR3X1_6 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_1_NAND3X1_220 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_42_DFFSR_49 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_31_DFFSR_89 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_8_DFFPOSX1_2 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_3_INVX1_83 INVX1_39/gnd DFFSR_54/S FILL
XNAND2X1_130 BUFX2_52/Y INVX1_169/A DFFSR_34/gnd OAI21X1_99/C DFFSR_34/S NAND2X1
XFILL_2_NOR2X1_66 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_50_DFFSR_105 INVX1_1/gnd DFFSR_53/S FILL
XFILL_7_DFFPOSX1_5 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_8_AOI21X1_22 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_43_5_0 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_6_DFFPOSX1_8 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_40_DFFSR_108 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_15_DFFSR_39 INVX1_3/gnd DFFSR_79/S FILL
XFILL_7_AOI21X1_25 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_2_NAND3X1_154 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_3_DFFSR_184 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_2_BUFX2_74 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_30_DFFSR_111 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_6_AOI21X1_28 AND2X2_38/B DFFSR_23/S FILL
XFILL_44_DFFSR_215 DFFSR_34/gnd DFFSR_1/S FILL
XDFFPOSX1_8 NOR3X1_3/A CLKBUF1_46/Y DFFPOSX1_8/D OR2X2_4/gnd DFFSR_32/S DFFPOSX1
XFILL_7_DFFPOSX1_28 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_20_DFFSR_114 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_5_AOI21X1_31 INVX1_39/gnd DFFSR_34/S FILL
XFILL_34_DFFSR_218 BUFX2_98/A DFFSR_32/S FILL
XFILL_10_DFFSR_117 BUFX2_77/gnd DFFSR_98/S FILL
XAOI21X1_28 AOI21X1_28/A AOI21X1_28/B AOI21X1_28/C AND2X2_38/B OAI21X1_73/B DFFSR_23/S
+ AOI21X1
XFILL_3_NAND2X1_5 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_24_DFFSR_221 AND2X2_38/B DFFSR_59/S FILL
XFILL_4_AOI21X1_34 INVX1_39/gnd DFFSR_34/S FILL
XFILL_50_DFFSR_56 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_39_DFFSR_96 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_3_AOI21X1_37 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_14_DFFSR_224 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_16_DFFPOSX1_47 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_2_AOI21X1_40 INVX1_39/gnd DFFSR_54/S FILL
XFILL_0_AND2X2_5 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_5_NAND2X1_124 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_6_DFFSR_53 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_6_DFFSR_111 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_12_DFFSR_86 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_1_AOI21X1_43 INVX1_3/gnd DFFSR_79/S FILL
XFILL_23_DFFSR_46 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_3_OAI22X1_4 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_47_DFFSR_142 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_0_AOI21X1_46 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_37_DFFSR_145 BUFX2_72/gnd DFFSR_201/S FILL
XBUFX2_31 BUFX2_34/A DFFSR_46/gnd BUFX2_31/Y DFFSR_54/S BUFX2
XFILL_0_DFFSR_221 AND2X2_38/B DFFSR_59/S FILL
XFILL_27_DFFSR_148 INVX1_67/gnd DFFSR_175/S FILL
XFILL_3_OAI21X1_106 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_26_DFFPOSX1_36 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_41_DFFSR_252 AND2X2_38/B DFFSR_23/S FILL
XFILL_3_INVX1_195 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_17_DFFSR_151 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_48_3 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_31_DFFSR_255 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_8_OAI21X1_70 INVX1_3/gnd DFFSR_23/S FILL
XFILL_1_NAND3X1_184 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_21_DFFSR_258 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_6_NAND2X1_91 INVX1_39/gnd DFFSR_54/S FILL
XFILL_7_OAI21X1_73 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_53_0_0 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_20_DFFSR_93 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_3_INVX1_47 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_42_DFFSR_13 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_31_DFFSR_53 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_2_NOR2X1_30 INVX1_3/gnd DFFSR_23/S FILL
XFILL_5_NAND2X1_94 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_6_OAI21X1_76 INVX1_1/gnd DFFSR_53/S FILL
XFILL_11_DFFSR_261 BUFX2_77/gnd DFFSR_98/S FILL
XNAND2X1_91 INVX1_162/Y NAND2X1_90/Y INVX1_39/gnd NAND2X1_91/Y DFFSR_54/S NAND2X1
XFILL_5_OAI21X1_79 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_4_NAND2X1_97 INVX1_1/gnd DFFSR_97/S FILL
XFILL_51_2_1 DFFSR_4/gnd DFFSR_98/S FILL
XOAI21X1_76 INVX1_166/Y XNOR2X1_3/A AOI22X1_26/A INVX1_1/gnd XOR2X1_6/A DFFSR_53/S
+ OAI21X1
XFILL_3_DFFSR_148 INVX1_67/gnd DFFSR_175/S FILL
XFILL_2_NAND3X1_118 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_4_OAI21X1_82 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_2_BUFX2_38 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_44_DFFSR_179 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_3_OAI21X1_85 INVX1_39/gnd DFFSR_54/S FILL
XFILL_7_DFFSR_255 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_4_NAND2X1_154 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_49_4_2 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_34_DFFSR_182 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_2_OAI21X1_88 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_21_DFFSR_4 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_24_DFFSR_185 INVX1_39/gnd DFFSR_54/S FILL
XFILL_0_INVX1_94 INVX1_67/gnd DFFSR_201/S FILL
XFILL_39_DFFSR_60 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_50_DFFSR_20 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_1_OAI21X1_91 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_14_DFFSR_188 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_0_OAI21X1_94 INVX1_67/gnd DFFSR_175/S FILL
XFILL_16_DFFPOSX1_11 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_6_DFFSR_17 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_23_DFFSR_10 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_12_DFFSR_50 BUFX2_77/gnd DFFSR_5/S FILL
XBUFX2_9 BUFX2_7/A AND2X2_38/B BUFX2_9/Y DFFSR_59/S BUFX2
XFILL_5_BUFX2_5 AND2X2_38/B DFFSR_59/S FILL
XFILL_47_DFFSR_106 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_0_NAND3X1_214 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_0_AOI21X1_10 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_37_DFFSR_109 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_17_3_0 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_0_DFFSR_185 INVX1_39/gnd DFFSR_54/S FILL
XFILL_27_DFFSR_112 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_41_DFFSR_216 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_3_INVX1_159 INVX1_3/gnd DFFSR_79/S FILL
XFILL_6_AND2X2_26 INVX1_1/gnd DFFSR_97/S FILL
XFILL_47_DFFSR_67 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_17_DFFSR_115 INVX1_1/gnd DFFSR_97/S FILL
XFILL_31_DFFSR_219 INVX1_67/gnd DFFSR_175/S FILL
XFILL_8_OAI21X1_34 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_1_NAND3X1_148 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_15_5_1 INVX1_39/gnd DFFSR_34/S FILL
XFILL_0_NAND2X1_6 BUFX2_98/A DFFSR_32/S FILL
XFILL_21_DFFSR_222 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_7_OAI21X1_37 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_6_NAND2X1_55 INVX1_39/gnd DFFSR_34/S FILL
XFILL_31_DFFSR_17 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_3_DFFSR_64 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_3_INVX1_11 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_20_DFFSR_57 BUFX2_79/A DFFSR_6/S FILL
XFILL_6_DFFPOSX1_22 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_5_NAND2X1_58 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_6_OAI21X1_40 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_11_DFFSR_225 INVX1_67/gnd DFFSR_175/S FILL
XNAND2X1_55 INVX1_62/A NAND2X1_55/B INVX1_39/gnd NAND2X1_55/Y DFFSR_34/S NAND2X1
XFILL_4_NAND2X1_61 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_5_OAI21X1_43 BUFX2_7/gnd DFFSR_151/S FILL
XOAI21X1_40 INVX1_143/A OAI21X1_40/B AOI22X1_20/A DFFSR_34/gnd AOI21X1_13/C DFFSR_1/S
+ OAI21X1
XFILL_3_DFFSR_112 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_4_OAI21X1_46 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_3_NAND2X1_64 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_0_OAI22X1_5 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_44_DFFSR_143 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_15_DFFPOSX1_41 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_2_NAND2X1_67 AND2X2_38/B DFFSR_59/S FILL
XFILL_3_OAI21X1_49 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_7_DFFSR_219 INVX1_67/gnd DFFSR_175/S FILL
XFILL_34_DFFSR_146 BUFX2_79/A DFFSR_7/S FILL
XFILL_4_NAND2X1_118 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_1_NAND2X1_70 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_2_OAI21X1_52 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_48_DFFSR_250 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_24_DFFSR_149 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_0_NAND2X1_73 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_39_DFFSR_24 BUFX2_98/A DFFSR_6/S FILL
XFILL_0_INVX1_58 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_10_AOI22X1_21 AND2X2_38/B DFFSR_59/S FILL
XFILL_0_INVX1_196 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_38_DFFSR_253 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_1_OAI21X1_55 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_28_DFFSR_64 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_14_DFFSR_152 INVX1_1/gnd DFFSR_53/S FILL
XFILL_28_DFFSR_256 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_0_OAI21X1_58 INVX1_39/gnd DFFSR_54/S FILL
XFILL_2_OAI21X1_100 INVX1_3/gnd DFFSR_79/S FILL
XFILL_25_DFFPOSX1_30 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_18_DFFSR_259 BUFX2_79/A DFFSR_6/S FILL
XFILL_9_AOI22X1_24 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_12_DFFSR_14 INVX1_1/gnd DFFSR_53/S FILL
XFILL_0_NAND3X1_178 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_8_AOI22X1_27 OR2X2_6/gnd DFFSR_92/S FILL
XNOR2X1_2 NOR3X1_1/A INVX1_3/Y INVX1_1/gnd NOR2X1_2/Y DFFSR_97/S NOR2X1
XFILL_0_DFFSR_149 BUFX2_72/gnd DFFSR_276/S FILL
XDFFSR_259 DFFSR_3/D DFFSR_3/CLK DFFSR_257/R DFFSR_6/S DFFSR_259/D BUFX2_79/A DFFSR_6/S
+ DFFSR
XFILL_25_0_1 AND2X2_38/B DFFSR_23/S FILL
XFILL_3_INVX1_123 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_41_DFFSR_180 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_47_DFFSR_31 BUFX2_79/A DFFSR_6/S FILL
XFILL_36_DFFSR_71 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_4_DFFSR_256 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_31_DFFSR_183 INVX1_67/gnd DFFSR_175/S FILL
XFILL_1_NAND3X1_112 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_23_2_2 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_6_NAND2X1_19 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_21_DFFSR_186 BUFX2_99/A DFFSR_92/S FILL
XFILL_3_DFFSR_28 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_20_DFFSR_21 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_3_NAND2X1_148 INVX1_67/gnd DFFSR_175/S FILL
XFILL_5_1_1 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_5_NAND2X1_22 BUFX2_99/A DFFSR_7/S FILL
XFILL_11_DFFSR_189 BUFX2_8/gnd DFFSR_51/S FILL
XNAND2X1_19 DFFSR_109/Q NOR2X1_5/Y DFFSR_8/gnd OAI21X1_5/C DFFSR_8/S NAND2X1
XFILL_4_NAND2X1_25 BUFX2_99/A DFFSR_7/S FILL
XFILL_6_NOR2X1_65 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_2_NOR2X1_9 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_3_3_2 INVX1_67/gnd DFFSR_175/S FILL
XFILL_9_DFFSR_3 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_4_OAI21X1_10 BUFX2_79/A DFFSR_7/S FILL
XFILL_3_NAND2X1_28 AND2X2_38/B DFFSR_59/S FILL
XDFFPOSX1_22 BUFX2_53/A CLKBUF1_49/Y NOR2X1_74/Y DFFSR_1/gnd DFFSR_81/S DFFPOSX1
XFILL_44_DFFSR_107 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_2_NAND2X1_31 INVX1_3/gnd DFFSR_23/S FILL
XFILL_3_OAI21X1_13 INVX1_39/gnd DFFSR_54/S FILL
XFILL_7_DFFSR_183 INVX1_67/gnd DFFSR_175/S FILL
XFILL_44_DFFSR_78 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_34_DFFSR_110 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_2_OAI21X1_16 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_1_NAND2X1_34 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_48_DFFSR_214 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_24_DFFSR_113 BUFX2_99/A DFFSR_92/S FILL
XFILL_8_NAND3X1_90 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_0_NAND2X1_37 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_1_OAI21X1_19 BUFX2_98/A DFFSR_32/S FILL
XFILL_38_DFFSR_217 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_0_INVX1_22 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_0_INVX1_160 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_0_DFFSR_75 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_28_DFFSR_28 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_17_DFFSR_68 BUFX2_98/A DFFSR_6/S FILL
XFILL_3_AND2X2_27 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_14_DFFSR_116 INVX1_3/gnd DFFSR_23/S FILL
XFILL_7_NAND3X1_93 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_28_DFFSR_220 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_0_OAI21X1_22 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_11_OAI22X1_9 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_6_NAND3X1_96 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_7_OR2X2_3 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_50_5_0 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_18_DFFSR_223 INVX1_39/gnd DFFSR_34/S FILL
XFILL_5_NAND3X1_99 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_0_NAND3X1_142 INVX1_67/gnd DFFSR_175/S FILL
XFILL_4_XOR2X1_5 OR2X2_6/gnd DFFSR_92/S FILL
XNAND3X1_96 NOR2X1_44/Y NOR2X1_45/Y NOR2X1_46/Y DFFSR_34/gnd INVX1_215/A DFFSR_1/S
+ NAND3X1
XFILL_33_DFFSR_7 BUFX2_79/A DFFSR_7/S FILL
XFILL_7_OAI22X1_3 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_5_DFFPOSX1_16 INVX1_67/gnd DFFSR_175/S FILL
XFILL_0_DFFSR_113 BUFX2_99/A DFFSR_92/S FILL
XFILL_2_NAND2X1_178 INVX1_1/gnd DFFSR_53/S FILL
XDFFSR_223 DFFSR_231/D CLKBUF1_29/Y BUFX2_66/Y DFFSR_34/S INVX1_106/A INVX1_39/gnd
+ DFFSR_34/S DFFSR
XFILL_41_DFFSR_144 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_36_DFFSR_35 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_8_DFFSR_82 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_25_DFFSR_75 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_4_DFFSR_220 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_31_DFFSR_147 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_45_DFFSR_251 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_21_DFFSR_150 AND2X2_38/B DFFSR_23/S FILL
XFILL_35_DFFSR_254 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_14_DFFPOSX1_35 INVX1_39/gnd DFFSR_54/S FILL
XFILL_3_NAND2X1_112 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_11_DFFSR_153 INVX1_67/gnd DFFSR_201/S FILL
XFILL_25_DFFSR_257 INVX1_39/gnd DFFSR_34/S FILL
XFILL_6_NOR2X1_29 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_15_DFFSR_260 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_0_NOR3X1_6 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_1_AOI22X1_12 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_10_OAI22X1_33 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_0_AOI22X1_15 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_33_DFFSR_82 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_44_DFFSR_42 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_7_DFFSR_147 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_24_DFFPOSX1_24 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_9_NAND3X1_51 BUFX2_99/A DFFSR_7/S FILL
XFILL_48_DFFSR_178 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_8_NAND3X1_54 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_9_OAI22X1_36 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_8_NAND3X1_227 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_0_DFFSR_39 INVX1_3/gnd DFFSR_79/S FILL
XFILL_38_DFFSR_181 INVX1_3/gnd DFFSR_79/S FILL
XFILL_0_INVX1_124 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_17_DFFSR_32 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_4_BUFX2_67 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_7_NAND3X1_57 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_8_OAI22X1_39 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_1_DFFSR_257 INVX1_39/gnd DFFSR_34/S FILL
XFILL_28_DFFSR_184 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_4_DFFPOSX1_46 INVX1_39/gnd DFFSR_34/S FILL
XFILL_6_NAND3X1_60 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_7_OAI22X1_42 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_18_DFFSR_187 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_6_OAI22X1_45 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_5_NAND3X1_63 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_0_NAND3X1_106 INVX1_3/gnd DFFSR_23/S FILL
XFILL_10_XOR2X1_2 OR2X2_2/gnd DFFSR_175/S FILL
XNAND3X1_60 NAND2X1_26/Y NAND3X1_60/B AND2X2_13/Y DFFSR_8/gnd NOR2X1_29/A DFFSR_8/S
+ NAND3X1
XFILL_4_NAND3X1_66 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_9_NAND3X1_161 AND2X2_38/B DFFSR_23/S FILL
XFILL_5_OAI22X1_48 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_41_DFFSR_89 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_3_NOR2X1_66 DFFSR_46/gnd DFFSR_62/S FILL
XOAI22X1_45 INVX1_108/Y OAI22X1_45/B INVX1_109/Y OAI22X1_45/D BUFX2_72/gnd NOR2X1_54/A
+ DFFSR_276/S OAI22X1
XFILL_51_DFFSR_105 INVX1_1/gnd DFFSR_53/S FILL
XFILL_3_NAND3X1_69 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_4_OAI22X1_51 INVX1_39/gnd DFFSR_54/S FILL
XFILL_2_NAND2X1_142 INVX1_67/gnd DFFSR_175/S FILL
XDFFSR_187 INVX1_77/A CLKBUF1_29/Y BUFX2_66/Y DFFSR_81/S DFFSR_187/D DFFSR_1/gnd DFFSR_81/S
+ DFFSR
XFILL_41_DFFSR_108 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_2_NAND3X1_72 INVX1_39/gnd DFFSR_34/S FILL
XFILL_25_DFFSR_39 INVX1_3/gnd DFFSR_79/S FILL
XFILL_8_DFFSR_46 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_14_DFFSR_79 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_4_DFFSR_184 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_31_DFFSR_111 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_1_NAND3X1_75 BUFX2_79/A DFFSR_7/S FILL
XFILL_45_DFFSR_215 DFFSR_34/gnd DFFSR_1/S FILL
XNAND2X1_8 INVX1_3/A NOR3X1_1/A INVX1_1/gnd NOR3X1_2/C DFFSR_53/S NAND2X1
XFILL_21_DFFSR_114 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_0_NAND3X1_78 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_35_DFFSR_218 BUFX2_98/A DFFSR_32/S FILL
XFILL_0_AND2X2_28 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_4_NAND2X1_5 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_11_DFFSR_117 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_25_DFFSR_221 AND2X2_38/B DFFSR_59/S FILL
XFILL_49_DFFSR_96 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_20_DFFSR_1 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_15_DFFSR_224 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_24_3_0 AND2X2_38/B DFFSR_59/S FILL
XOAI22X1_7 INVX1_17/Y OAI22X1_7/B INVX1_18/Y OAI22X1_7/D AND2X2_38/B OAI22X1_7/Y DFFSR_59/S
+ OAI22X1
XINVX1_80 INVX1_80/A DFFSR_1/gnd INVX1_80/Y DFFSR_81/S INVX1
XFILL_7_DFFSR_111 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_5_DFFSR_93 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_22_DFFSR_86 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_33_DFFSR_46 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_4_OAI22X1_4 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_48_DFFSR_142 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_22_5_1 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_8_NAND3X1_18 BUFX2_79/A DFFSR_7/S FILL
XFILL_4_BUFX2_2 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_38_DFFSR_145 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_8_NAND3X1_191 BUFX2_7/gnd DFFSR_151/S FILL
XINVX1_198 BUFX2_38/Y DFFSR_34/gnd DFFSR_266/R DFFSR_1/S INVX1
XFILL_4_4_0 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_7_NAND3X1_21 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_1_DFFSR_221 AND2X2_38/B DFFSR_59/S FILL
XFILL_4_BUFX2_31 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_4_DFFPOSX1_10 INVX1_67/gnd DFFSR_201/S FILL
XFILL_28_DFFSR_148 INVX1_67/gnd DFFSR_175/S FILL
XFILL_42_DFFSR_252 AND2X2_38/B DFFSR_23/S FILL
XFILL_1_NAND2X1_172 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_6_NAND3X1_24 INVX1_1/gnd DFFSR_97/S FILL
XFILL_18_DFFSR_151 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_32_DFFSR_255 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_2_6_1 INVX1_67/gnd DFFSR_201/S FILL
XFILL_5_NAND3X1_27 OR2X2_4/gnd DFFSR_3/S FILL
XNAND3X1_24 NOR2X1_12/Y NOR2X1_13/Y NOR2X1_14/Y INVX1_1/gnd XOR2X1_10/A DFFSR_97/S
+ NAND3X1
XFILL_22_DFFSR_258 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_4_NAND3X1_30 BUFX2_79/A DFFSR_6/S FILL
XFILL_2_INVX1_87 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_5_OAI22X1_12 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_41_DFFSR_53 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_30_DFFSR_93 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_3_NOR2X1_30 INVX1_3/gnd DFFSR_23/S FILL
XFILL_13_DFFPOSX1_29 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_12_DFFSR_261 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_4_OAI22X1_15 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_3_NAND3X1_33 DFFSR_8/gnd DFFSR_8/S FILL
XDFFSR_151 DFFSR_167/D CLKBUF1_14/Y BUFX2_64/Y DFFSR_151/S DFFSR_151/D XOR2X1_1/gnd
+ DFFSR_151/S DFFSR
XFILL_2_NAND2X1_106 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_3_OAI22X1_18 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_2_NAND3X1_36 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_8_DFFSR_10 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_4_DFFSR_148 INVX1_67/gnd DFFSR_175/S FILL
XFILL_14_DFFSR_43 BUFX2_98/A DFFSR_6/S FILL
XFILL_1_BUFX2_78 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_1_NAND3X1_39 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_2_OAI22X1_21 BUFX2_98/A DFFSR_32/S FILL
XFILL_45_DFFSR_179 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_8_DFFSR_255 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_1_OAI22X1_24 BUFX2_98/A DFFSR_32/S FILL
XFILL_0_NAND3X1_42 BUFX2_79/A DFFSR_6/S FILL
XFILL_35_DFFSR_182 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_23_DFFPOSX1_18 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_0_OAI22X1_27 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_25_DFFSR_185 INVX1_39/gnd DFFSR_54/S FILL
XFILL_49_DFFSR_60 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_7_NAND3X1_221 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_15_DFFSR_188 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_3_DFFPOSX1_40 OR2X2_1/gnd DFFSR_59/S FILL
XINVX1_44 INVX1_44/A OR2X2_4/gnd INVX1_44/Y DFFSR_3/S INVX1
XFILL_32_0_1 INVX1_1/gnd DFFSR_97/S FILL
XDFFSR_97 DFFSR_97/Q DFFSR_83/CLK DFFSR_73/R DFFSR_97/S DFFSR_89/Q INVX1_1/gnd DFFSR_97/S
+ DFFSR
XFILL_33_DFFSR_10 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_22_DFFSR_50 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_11_DFFSR_90 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_5_DFFSR_57 BUFX2_79/A DFFSR_6/S FILL
XFILL_0_NOR2X1_67 INVX1_67/gnd DFFSR_175/S FILL
XFILL_48_DFFSR_106 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_8_NAND3X1_155 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_38_DFFSR_109 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_30_2_2 XOR2X1_4/gnd DFFSR_91/S FILL
XINVX1_162 INVX1_162/A INVX1_39/gnd INVX1_162/Y DFFSR_34/S INVX1
XFILL_1_DFFSR_185 INVX1_39/gnd DFFSR_54/S FILL
XFILL_28_DFFSR_112 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_1_NAND2X1_136 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_42_DFFSR_216 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_4_INVX1_159 INVX1_3/gnd DFFSR_79/S FILL
XFILL_7_AND2X2_26 INVX1_1/gnd DFFSR_97/S FILL
XFILL_18_DFFSR_115 INVX1_1/gnd DFFSR_97/S FILL
XFILL_32_DFFSR_219 INVX1_67/gnd DFFSR_175/S FILL
XFILL_1_NAND2X1_6 BUFX2_98/A DFFSR_32/S FILL
XFILL_22_DFFSR_222 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_41_DFFSR_17 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_2_INVX1_51 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_30_DFFSR_57 BUFX2_79/A DFFSR_6/S FILL
XFILL_19_DFFSR_97 INVX1_1/gnd DFFSR_97/S FILL
XFILL_12_DFFSR_225 INVX1_67/gnd DFFSR_175/S FILL
XDFFSR_115 INVX1_23/A CLKBUF1_27/Y BUFX2_49/Y DFFSR_97/S DFFSR_115/D INVX1_1/gnd DFFSR_97/S
+ DFFSR
XFILL_22_DFFPOSX1_48 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_4_DFFSR_112 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_1_BUFX2_42 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_1_OAI22X1_5 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_45_DFFSR_143 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_8_DFFSR_219 INVX1_67/gnd DFFSR_175/S FILL
XFILL_35_DFFSR_146 BUFX2_79/A DFFSR_7/S FILL
XFILL_49_DFFSR_250 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_11_DFFSR_8 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_25_DFFSR_149 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_39_DFFSR_253 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_38_DFFSR_64 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_49_DFFSR_24 BUFX2_98/A DFFSR_6/S FILL
XFILL_1_INVX1_196 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_7_NAND3X1_185 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_15_DFFSR_152 INVX1_1/gnd DFFSR_53/S FILL
XFILL_29_DFFSR_256 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_0_NAND2X1_166 BUFX2_8/gnd DFFSR_81/S FILL
XDFFSR_61 INVX1_32/A DFFSR_57/CLK DFFSR_35/R DFFSR_8/S DFFSR_61/D DFFSR_28/gnd DFFSR_8/S
+ DFFSR
XFILL_5_DFFSR_21 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_19_DFFSR_259 BUFX2_79/A DFFSR_6/S FILL
XFILL_22_DFFSR_14 INVX1_1/gnd DFFSR_53/S FILL
XFILL_11_DFFSR_54 INVX1_39/gnd DFFSR_54/S FILL
XFILL_0_NOR2X1_31 INVX1_39/gnd DFFSR_54/S FILL
XINVX1_126 NOR3X1_4/A INVX1_3/gnd INVX1_126/Y DFFSR_23/S INVX1
XFILL_8_NAND3X1_119 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_4_NOR2X1_2 INVX1_1/gnd DFFSR_97/S FILL
XFILL_1_DFFSR_149 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_12_DFFPOSX1_23 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_32_DFFSR_4 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_42_DFFSR_180 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_1_NAND2X1_100 INVX1_39/gnd DFFSR_54/S FILL
XFILL_46_DFFSR_71 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_5_DFFSR_256 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_32_DFFSR_183 INVX1_67/gnd DFFSR_175/S FILL
XFILL_22_DFFSR_186 BUFX2_99/A DFFSR_92/S FILL
XFILL_30_DFFSR_21 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_2_INVX1_15 BUFX2_98/A DFFSR_32/S FILL
XFILL_2_DFFSR_68 BUFX2_98/A DFFSR_6/S FILL
XFILL_19_DFFSR_61 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_6_BUFX2_96 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_12_DFFSR_189 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_22_DFFPOSX1_12 AND2X2_38/B DFFSR_23/S FILL
XFILL_6_NAND3X1_215 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_45_DFFSR_107 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_2_DFFPOSX1_34 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_8_DFFSR_183 INVX1_67/gnd DFFSR_175/S FILL
XFILL_35_DFFSR_110 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_49_DFFSR_214 BUFX2_72/gnd DFFSR_276/S FILL
XAND2X2_30 NOR2X1_67/Y AND2X2_30/B OR2X2_2/gnd AND2X2_30/Y DFFSR_175/S AND2X2
XFILL_25_DFFSR_113 BUFX2_99/A DFFSR_92/S FILL
XFILL_39_DFFSR_217 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_38_DFFSR_28 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_27_DFFSR_68 BUFX2_98/A DFFSR_6/S FILL
XFILL_1_INVX1_160 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_4_AND2X2_27 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_15_DFFSR_116 INVX1_3/gnd DFFSR_23/S FILL
XFILL_7_NAND3X1_149 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_29_DFFSR_220 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_0_NAND2X1_130 DFFSR_34/gnd DFFSR_34/S FILL
XDFFSR_25 INVX1_8/A CLKBUF1_7/Y DFFSR_3/R DFFSR_3/S DFFSR_1/Q OR2X2_4/gnd DFFSR_3/S
+ DFFSR
XFILL_19_DFFSR_223 INVX1_39/gnd DFFSR_34/S FILL
XFILL_11_DFFSR_18 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_8_OAI22X1_3 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_17_2 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_1_DFFSR_113 BUFX2_99/A DFFSR_92/S FILL
XFILL_21_DFFPOSX1_42 INVX1_39/gnd DFFSR_34/S FILL
XFILL_42_DFFSR_144 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_46_DFFSR_35 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_35_DFFSR_75 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_5_DFFSR_220 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_32_DFFSR_147 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_46_DFFSR_251 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_5_NAND3X1_245 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_22_DFFSR_150 AND2X2_38/B DFFSR_23/S FILL
XFILL_31_3_0 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_2_DFFSR_32 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_36_DFFSR_254 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_19_DFFSR_25 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_12_DFFSR_153 INVX1_67/gnd DFFSR_201/S FILL
XFILL_6_BUFX2_60 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_26_DFFSR_257 INVX1_39/gnd DFFSR_34/S FILL
XFILL_8_OAI21X1_101 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_29_5_1 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_16_DFFSR_260 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_20_CLKBUF1_15 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_6_NAND3X1_179 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_43_DFFSR_82 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_19_CLKBUF1_18 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_8_DFFSR_147 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_18_CLKBUF1_21 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_49_DFFSR_178 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_9_6_1 XOR2X1_1/gnd DFFSR_208/S FILL
XNAND3X1_215 NAND3X1_215/A NAND3X1_215/B OAI21X1_59/Y DFFSR_62/gnd NAND3X1_215/Y DFFSR_62/S
+ NAND3X1
XFILL_17_CLKBUF1_24 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_39_DFFSR_181 INVX1_3/gnd DFFSR_79/S FILL
XFILL_1_INVX1_124 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_16_DFFSR_72 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_27_DFFSR_32 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_2_DFFSR_257 INVX1_39/gnd DFFSR_34/S FILL
XFILL_7_NAND3X1_113 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_16_CLKBUF1_27 INVX1_1/gnd DFFSR_97/S FILL
XFILL_29_DFFSR_184 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_11_DFFPOSX1_17 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_15_CLKBUF1_30 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_19_DFFSR_187 DFFSR_1/gnd DFFSR_81/S FILL
XNOR2X1_69 INVX1_134/Y NOR2X1_69/B OR2X2_6/gnd NOR2X1_69/Y DFFSR_92/S NOR2X1
XFILL_14_CLKBUF1_33 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_3_XOR2X1_9 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_51_DFFSR_89 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_13_CLKBUF1_36 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_4_NOR2X1_66 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_12_CLKBUF1_39 INVX1_1/gnd DFFSR_53/S FILL
XFILL_42_DFFSR_108 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_7_DFFSR_86 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_11_CLKBUF1_42 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_24_DFFSR_79 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_35_DFFSR_39 INVX1_3/gnd DFFSR_79/S FILL
XFILL_5_DFFSR_184 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_32_DFFSR_111 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_10_CLKBUF1_45 BUFX2_79/A DFFSR_7/S FILL
XFILL_46_DFFSR_215 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_5_NAND3X1_209 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_22_DFFSR_114 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_1_DFFPOSX1_28 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_36_DFFSR_218 BUFX2_98/A DFFSR_32/S FILL
XFILL_39_0_1 BUFX2_79/A DFFSR_6/S FILL
XFILL_1_AND2X2_28 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_6_BUFX2_24 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_5_NAND2X1_5 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_12_DFFSR_117 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_9_CLKBUF1_48 INVX1_3/gnd DFFSR_79/S FILL
XFILL_26_DFFSR_221 AND2X2_38/B DFFSR_59/S FILL
XFILL_16_DFFSR_224 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_44_DFFSR_7 BUFX2_79/A DFFSR_7/S FILL
XFILL_16_NOR3X1_3 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_37_2_2 BUFX2_99/A DFFSR_7/S FILL
XFILL_6_NAND3X1_143 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_10_DFFPOSX1_47 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_8_DFFSR_111 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_32_DFFSR_86 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_4_INVX1_80 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_43_DFFSR_46 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_5_OAI22X1_4 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_49_DFFSR_142 XOR2X1_1/gnd DFFSR_151/S FILL
XNAND3X1_179 INVX1_160/Y NAND3X1_176/B NAND3X1_176/C NOR3X1_6/gnd AOI21X1_27/B DFFSR_79/S
+ NAND3X1
XFILL_39_DFFSR_145 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_16_DFFSR_36 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_2_DFFSR_221 AND2X2_38/B DFFSR_59/S FILL
XFILL_29_DFFSR_148 INVX1_67/gnd DFFSR_175/S FILL
XFILL_3_BUFX2_71 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_39_2 BUFX2_79/A DFFSR_7/S FILL
XFILL_43_DFFSR_252 AND2X2_38/B DFFSR_23/S FILL
XFILL_20_DFFPOSX1_36 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_19_DFFSR_151 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_33_DFFSR_255 OR2X2_4/gnd DFFSR_32/S FILL
XNOR2X1_33 INVX1_62/A NOR3X1_3/A INVX1_3/gnd AND2X2_18/B DFFSR_23/S NOR2X1
XFILL_4_NAND3X1_239 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_23_DFFSR_258 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_40_DFFSR_93 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_4_NOR2X1_30 INVX1_3/gnd DFFSR_23/S FILL
XFILL_13_DFFSR_261 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_1_AND2X2_2 BUFX2_99/A DFFSR_7/S FILL
XFILL_7_DFFSR_50 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_24_DFFSR_43 BUFX2_98/A DFFSR_6/S FILL
XFILL_13_DFFSR_83 INVX1_3/gnd DFFSR_79/S FILL
XFILL_5_DFFSR_148 INVX1_67/gnd DFFSR_175/S FILL
XFILL_5_NAND3X1_173 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_46_DFFSR_179 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_9_DFFSR_255 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_36_DFFSR_182 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_9_CLKBUF1_12 AND2X2_38/B DFFSR_23/S FILL
XFILL_26_DFFSR_185 INVX1_39/gnd DFFSR_54/S FILL
XFILL_10_DFFSR_5 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_16_DFFSR_188 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_8_CLKBUF1_15 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_6_NAND3X1_107 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_7_CLKBUF1_18 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_10_DFFPOSX1_11 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_43_DFFSR_10 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_32_DFFSR_50 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_4_INVX1_44 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_4_DFFSR_97 INVX1_1/gnd DFFSR_97/S FILL
XFILL_21_DFFSR_90 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_1_NOR2X1_67 INVX1_67/gnd DFFSR_175/S FILL
XFILL_6_CLKBUF1_21 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_49_DFFSR_106 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_5_CLKBUF1_24 DFFSR_4/gnd DFFSR_98/S FILL
XNAND3X1_143 AOI22X1_19/C INVX1_144/Y OAI21X1_38/C BUFX2_8/gnd AOI21X1_12/B DFFSR_51/S
+ NAND3X1
XFILL_39_DFFSR_109 DFFSR_4/gnd DFFSR_4/S FILL
XCLKBUF1_21 BUFX2_3/Y XOR2X1_1/gnd CLKBUF1_21/Y DFFSR_151/S CLKBUF1
XFILL_4_CLKBUF1_27 INVX1_1/gnd DFFSR_97/S FILL
XOR2X2_1 OR2X2_1/A OR2X2_1/B OR2X2_1/gnd OR2X2_1/Y DFFSR_59/S OR2X2
XFILL_2_DFFSR_185 INVX1_39/gnd DFFSR_54/S FILL
XFILL_29_DFFSR_112 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_3_BUFX2_35 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_43_DFFSR_216 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_3_CLKBUF1_30 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_8_AND2X2_26 INVX1_1/gnd DFFSR_97/S FILL
XFILL_19_DFFSR_115 INVX1_1/gnd DFFSR_97/S FILL
XFILL_33_DFFSR_219 INVX1_67/gnd DFFSR_175/S FILL
XFILL_2_CLKBUF1_33 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_31_DFFSR_1 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_2_NAND2X1_6 BUFX2_98/A DFFSR_32/S FILL
XFILL_23_DFFSR_222 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_4_NAND3X1_203 INVX1_1/gnd DFFSR_97/S FILL
XFILL_1_CLKBUF1_36 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_51_DFFSR_17 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_40_DFFSR_57 BUFX2_79/A DFFSR_6/S FILL
XFILL_29_DFFSR_97 INVX1_1/gnd DFFSR_97/S FILL
XFILL_1_INVX1_91 AND2X2_38/B DFFSR_23/S FILL
XFILL_13_DFFSR_225 INVX1_67/gnd DFFSR_175/S FILL
XFILL_0_CLKBUF1_39 INVX1_1/gnd DFFSR_53/S FILL
XFILL_0_DFFPOSX1_22 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_11_0_2 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_7_DFFSR_14 INVX1_1/gnd DFFSR_53/S FILL
XFILL_13_DFFSR_47 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_5_DFFSR_112 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_0_BUFX2_82 INVX1_1/gnd DFFSR_97/S FILL
XFILL_2_OAI22X1_5 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_46_DFFSR_143 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_5_NAND3X1_137 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_9_DFFSR_219 INVX1_67/gnd DFFSR_175/S FILL
XFILL_36_DFFSR_146 BUFX2_79/A DFFSR_7/S FILL
XFILL_50_DFFSR_250 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_26_DFFSR_149 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_40_DFFSR_253 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_48_DFFSR_64 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_2_INVX1_196 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_16_DFFSR_152 INVX1_1/gnd DFFSR_53/S FILL
XFILL_30_DFFSR_256 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_20_DFFSR_259 BUFX2_79/A DFFSR_6/S FILL
XFILL_4_DFFSR_61 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_32_DFFSR_14 INVX1_1/gnd DFFSR_53/S FILL
XFILL_19_DFFPOSX1_30 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_10_DFFSR_94 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_21_DFFSR_54 INVX1_39/gnd DFFSR_54/S FILL
XFILL_1_NOR2X1_31 INVX1_39/gnd DFFSR_54/S FILL
XFILL_10_DFFSR_262 BUFX2_98/A DFFSR_32/S FILL
XNAND3X1_107 BUFX2_95/A AND2X2_16/Y BUFX2_32/Y BUFX2_8/gnd AND2X2_24/A DFFSR_81/S
+ NAND3X1
XFILL_3_NAND3X1_233 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_38_3_0 BUFX2_79/A DFFSR_7/S FILL
XFILL_2_DFFSR_149 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_43_DFFSR_180 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_6_DFFSR_256 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_33_DFFSR_183 INVX1_67/gnd DFFSR_175/S FILL
XFILL_36_5_1 BUFX2_99/A DFFSR_92/S FILL
XFILL_23_DFFSR_186 BUFX2_99/A DFFSR_92/S FILL
XFILL_4_NAND3X1_167 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_29_DFFSR_61 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_1_INVX1_55 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_40_DFFSR_21 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_13_DFFSR_189 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_9_DFFPOSX1_41 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_13_DFFSR_11 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_0_BUFX2_46 BUFX2_98/A DFFSR_6/S FILL
XFILL_46_DFFSR_107 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_5_NAND3X1_101 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_9_DFFSR_183 INVX1_67/gnd DFFSR_175/S FILL
XFILL_36_DFFSR_110 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_50_DFFSR_214 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_26_DFFSR_113 BUFX2_99/A DFFSR_92/S FILL
XFILL_40_DFFSR_217 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_48_DFFSR_28 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_37_DFFSR_68 BUFX2_98/A DFFSR_6/S FILL
XFILL_2_INVX1_160 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_5_AND2X2_27 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_16_DFFSR_116 INVX1_3/gnd DFFSR_23/S FILL
XFILL_30_DFFSR_220 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_20_DFFSR_223 INVX1_39/gnd DFFSR_34/S FILL
XFILL_4_DFFSR_25 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_21_DFFSR_18 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_10_DFFSR_58 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_5_OAI21X1_119 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_10_DFFSR_226 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_3_NAND3X1_197 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_9_OAI22X1_3 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_3_NOR2X1_6 BUFX2_98/A DFFSR_6/S FILL
XFILL_2_DFFSR_113 BUFX2_99/A DFFSR_92/S FILL
XFILL_46_0_1 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_22_DFFSR_8 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_43_DFFSR_144 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_45_DFFSR_75 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_6_DFFSR_220 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_33_DFFSR_147 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_47_DFFSR_251 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_44_2_2 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_23_DFFSR_150 AND2X2_38/B DFFSR_23/S FILL
XFILL_4_NAND3X1_131 AND2X2_38/B DFFSR_59/S FILL
XFILL_1_INVX1_19 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_1_DFFSR_72 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_29_DFFSR_25 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_18_DFFSR_65 BUFX2_79/A DFFSR_7/S FILL
XFILL_37_DFFSR_254 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_13_DFFSR_153 INVX1_67/gnd DFFSR_201/S FILL
XFILL_6_BUFX2_9 AND2X2_38/B DFFSR_59/S FILL
XFILL_27_DFFSR_257 INVX1_39/gnd DFFSR_34/S FILL
XFILL_6_NAND2X1_167 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_17_DFFSR_260 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_0_BUFX2_10 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_5_XOR2X1_2 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_43_DFFSR_4 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_9_DFFSR_147 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_18_DFFPOSX1_24 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_20_DFFPOSX1_3 INVX1_39/gnd DFFSR_34/S FILL
XFILL_50_DFFSR_178 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_19_DFFPOSX1_6 AND2X2_38/B DFFSR_23/S FILL
XFILL_12_1_0 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_40_DFFSR_181 INVX1_3/gnd DFFSR_79/S FILL
XFILL_37_DFFSR_32 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_9_DFFSR_79 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_2_INVX1_124 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_26_DFFSR_72 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_2_NAND3X1_227 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_18_DFFPOSX1_9 INVX1_67/gnd DFFSR_201/S FILL
XFILL_3_DFFSR_257 INVX1_39/gnd DFFSR_34/S FILL
XFILL_30_DFFSR_184 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_10_3_1 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_20_DFFSR_187 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_10_DFFSR_22 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_10_DFFSR_190 INVX1_39/gnd DFFSR_34/S FILL
XFILL_3_NAND3X1_161 AND2X2_38/B DFFSR_23/S FILL
XFILL_5_NOR2X1_66 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_1_NOR3X1_3 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_43_DFFSR_108 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_8_DFFPOSX1_35 INVX1_39/gnd DFFSR_54/S FILL
XFILL_34_DFFSR_79 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_45_DFFSR_39 INVX1_3/gnd DFFSR_79/S FILL
XFILL_6_DFFSR_184 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_33_DFFSR_111 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_47_DFFSR_215 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_23_DFFSR_114 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_37_DFFSR_218 BUFX2_98/A DFFSR_32/S FILL
XFILL_18_DFFSR_29 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_1_DFFSR_36 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_2_AND2X2_28 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_6_NAND2X1_5 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_13_DFFSR_117 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_5_BUFX2_64 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_27_DFFSR_221 AND2X2_38/B DFFSR_59/S FILL
XFILL_6_NAND2X1_131 INVX1_3/gnd DFFSR_79/S FILL
XFILL_17_DFFSR_224 BUFX2_7/gnd DFFSR_151/S FILL
XXOR2X1_6 XOR2X1_6/A XOR2X1_5/Y BUFX2_99/A XOR2X1_6/Y DFFSR_7/S XOR2X1
XFILL_42_DFFSR_86 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_9_DFFSR_111 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_9_AOI21X1_56 NOR3X1_6/gnd DFFSR_79/S FILL
XNAND2X1_167 DFFSR_59/S NAND2X1_167/B OR2X2_1/gnd AOI21X1_59/B DFFSR_59/S NAND2X1
XFILL_6_OAI22X1_4 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_50_DFFSR_142 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_4_OAI21X1_113 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_8_AOI21X1_59 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_27_DFFPOSX1_43 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_40_DFFSR_145 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_9_DFFSR_43 BUFX2_98/A DFFSR_6/S FILL
XFILL_7_AOI21X1_62 INVX1_3/gnd DFFSR_23/S FILL
XFILL_2_NAND3X1_191 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_26_DFFSR_36 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_15_DFFSR_76 BUFX2_79/A DFFSR_7/S FILL
XFILL_3_DFFSR_221 AND2X2_38/B DFFSR_59/S FILL
XFILL_30_DFFSR_148 INVX1_67/gnd DFFSR_175/S FILL
XFILL_6_AOI21X1_65 INVX1_3/gnd DFFSR_23/S FILL
XFILL_44_DFFSR_252 AND2X2_38/B DFFSR_23/S FILL
XFILL_20_DFFSR_151 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_5_AOI21X1_68 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_34_DFFSR_255 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_18_0_2 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_10_DFFSR_154 BUFX2_99/A DFFSR_7/S FILL
XAOI21X1_65 AOI21X1_64/A XOR2X1_10/Y AND2X2_42/Y INVX1_3/gnd XOR2X1_12/A DFFSR_23/S
+ AOI21X1
XFILL_4_AOI21X1_71 BUFX2_99/A DFFSR_92/S FILL
XFILL_24_DFFSR_258 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_50_DFFSR_93 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_3_NAND3X1_125 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_5_NOR2X1_30 INVX1_3/gnd DFFSR_23/S FILL
XFILL_14_DFFSR_261 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_5_NAND2X1_161 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_6_DFFSR_90 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_34_DFFSR_43 BUFX2_98/A DFFSR_6/S FILL
XFILL_23_DFFSR_83 INVX1_3/gnd DFFSR_79/S FILL
XFILL_6_DFFSR_148 INVX1_67/gnd DFFSR_175/S FILL
XFILL_47_DFFSR_179 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_37_DFFSR_182 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_0_DFFSR_258 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_5_BUFX2_28 DFFSR_46/gnd DFFSR_62/S FILL
XBUFX2_68 BUFX2_60/A XOR2X1_1/gnd BUFX2_68/Y DFFSR_208/S BUFX2
XFILL_17_DFFPOSX1_18 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_27_DFFSR_185 INVX1_39/gnd DFFSR_54/S FILL
XFILL_17_DFFSR_188 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_1_NAND3X1_221 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_45_3_0 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_42_DFFSR_50 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_8_DFFPOSX1_3 INVX1_39/gnd DFFSR_34/S FILL
XFILL_3_INVX1_84 INVX1_39/gnd DFFSR_34/S FILL
XFILL_31_DFFSR_90 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_9_AOI21X1_20 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_2_NOR2X1_67 INVX1_67/gnd DFFSR_175/S FILL
XNAND2X1_131 BUFX2_55/Y INVX1_180/A INVX1_3/gnd NAND2X1_131/Y DFFSR_79/S NAND2X1
XFILL_50_DFFSR_106 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_7_DFFPOSX1_6 AND2X2_38/B DFFSR_23/S FILL
XFILL_8_AOI21X1_23 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_43_5_1 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_40_DFFSR_109 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_6_DFFPOSX1_9 INVX1_67/gnd DFFSR_201/S FILL
XFILL_7_AOI21X1_26 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_2_NAND3X1_155 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_15_DFFSR_40 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_3_DFFSR_185 INVX1_39/gnd DFFSR_54/S FILL
XFILL_2_BUFX2_75 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_30_DFFSR_112 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_44_DFFSR_216 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_6_AOI21X1_29 DFFSR_62/gnd DFFSR_208/S FILL
XDFFPOSX1_9 INVX1_62/A CLKBUF1_43/Y DFFPOSX1_9/D INVX1_67/gnd DFFSR_201/S DFFPOSX1
XFILL_9_AND2X2_26 INVX1_1/gnd DFFSR_97/S FILL
XFILL_7_DFFPOSX1_29 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_20_DFFSR_115 INVX1_1/gnd DFFSR_97/S FILL
XFILL_5_AOI21X1_32 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_34_DFFSR_219 INVX1_67/gnd DFFSR_175/S FILL
XFILL_10_DFFSR_118 OR2X2_3/gnd DFFSR_60/S FILL
XAOI21X1_29 AOI21X1_29/A AOI21X1_29/B OAI21X1_54/C DFFSR_62/gnd AOI21X1_29/Y DFFSR_208/S
+ AOI21X1
XFILL_3_NAND2X1_6 BUFX2_98/A DFFSR_32/S FILL
XFILL_4_AOI21X1_35 INVX1_39/gnd DFFSR_54/S FILL
XFILL_24_DFFSR_222 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_50_DFFSR_57 BUFX2_79/A DFFSR_6/S FILL
XFILL_39_DFFSR_97 INVX1_1/gnd DFFSR_97/S FILL
XFILL_3_AOI21X1_38 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_14_DFFSR_225 INVX1_67/gnd DFFSR_175/S FILL
XFILL_16_DFFPOSX1_48 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_2_AOI21X1_41 INVX1_39/gnd DFFSR_34/S FILL
XFILL_0_AND2X2_6 BUFX2_99/A DFFSR_7/S FILL
XFILL_5_NAND2X1_125 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_23_DFFSR_47 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_6_DFFSR_54 INVX1_39/gnd DFFSR_54/S FILL
XFILL_1_AOI21X1_44 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_12_DFFSR_87 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_6_DFFSR_112 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_3_OAI22X1_5 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_47_DFFSR_143 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_0_AOI21X1_47 INVX1_67/gnd DFFSR_175/S FILL
XFILL_37_DFFSR_146 BUFX2_79/A DFFSR_7/S FILL
XFILL_0_DFFSR_222 BUFX2_72/gnd DFFSR_201/S FILL
XBUFX2_32 BUFX2_34/A BUFX2_8/gnd BUFX2_32/Y DFFSR_51/S BUFX2
XFILL_27_DFFSR_149 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_3_OAI21X1_107 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_26_DFFPOSX1_37 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_3_INVX1_196 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_41_DFFSR_253 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_48_4 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_17_DFFSR_152 INVX1_1/gnd DFFSR_53/S FILL
XFILL_8_OAI21X1_71 INVX1_3/gnd DFFSR_79/S FILL
XFILL_1_NAND3X1_185 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_31_DFFSR_256 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_6_NAND2X1_92 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_21_DFFSR_259 BUFX2_79/A DFFSR_6/S FILL
XFILL_7_OAI21X1_74 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_3_INVX1_48 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_53_0_1 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_42_DFFSR_14 INVX1_1/gnd DFFSR_53/S FILL
XFILL_20_DFFSR_94 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_31_DFFSR_54 INVX1_39/gnd DFFSR_54/S FILL
XFILL_2_NOR2X1_31 INVX1_39/gnd DFFSR_54/S FILL
XFILL_6_OAI21X1_77 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_11_DFFSR_262 BUFX2_98/A DFFSR_32/S FILL
XFILL_5_NAND2X1_95 XOR2X1_4/gnd DFFSR_91/S FILL
XNAND2X1_92 INVX1_145/A AND2X2_35/B NOR3X1_6/gnd XOR2X1_4/A DFFSR_79/S NAND2X1
XFILL_5_OAI21X1_80 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_4_NAND2X1_98 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_51_2_2 DFFSR_4/gnd DFFSR_98/S FILL
XOAI21X1_77 INVX1_175/Y INVX1_161/Y XNOR2X1_2/Y DFFSR_8/gnd OAI21X1_77/Y DFFSR_8/S
+ OAI21X1
XFILL_2_NAND3X1_119 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_3_DFFSR_149 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_4_OAI21X1_83 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_2_BUFX2_39 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_44_DFFSR_180 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_3_OAI21X1_86 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_7_DFFSR_256 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_4_NAND2X1_155 BUFX2_79/A DFFSR_7/S FILL
XFILL_34_DFFSR_183 INVX1_67/gnd DFFSR_175/S FILL
XFILL_2_OAI21X1_89 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_21_DFFSR_5 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_24_DFFSR_186 BUFX2_99/A DFFSR_92/S FILL
XFILL_1_OAI21X1_92 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_0_INVX1_95 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_39_DFFSR_61 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_50_DFFSR_21 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_14_DFFSR_189 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_0_OAI21X1_95 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_16_DFFPOSX1_12 AND2X2_38/B DFFSR_23/S FILL
XFILL_6_DFFSR_18 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_19_1_0 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_23_DFFSR_11 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_5_BUFX2_6 BUFX2_79/A DFFSR_6/S FILL
XFILL_12_DFFSR_51 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_47_DFFSR_107 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_0_NAND3X1_215 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_0_AOI21X1_11 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_37_DFFSR_110 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_17_3_1 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_51_DFFSR_214 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_0_DFFSR_186 BUFX2_99/A DFFSR_92/S FILL
XFILL_27_DFFSR_113 BUFX2_99/A DFFSR_92/S FILL
XFILL_41_DFFSR_217 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_9_OAI21X1_32 AND2X2_38/B DFFSR_59/S FILL
XFILL_42_DFFSR_1 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_47_DFFSR_68 BUFX2_98/A DFFSR_6/S FILL
XFILL_3_INVX1_160 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_6_AND2X2_27 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_17_DFFSR_116 INVX1_3/gnd DFFSR_23/S FILL
XFILL_8_OAI21X1_35 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_15_5_2 INVX1_39/gnd DFFSR_34/S FILL
XFILL_31_DFFSR_220 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_1_NAND3X1_149 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_0_NAND2X1_7 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_6_NAND2X1_56 AND2X2_38/B DFFSR_59/S FILL
XFILL_7_OAI21X1_38 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_21_DFFSR_223 INVX1_39/gnd DFFSR_34/S FILL
XFILL_3_INVX1_12 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_3_DFFSR_65 BUFX2_79/A DFFSR_7/S FILL
XFILL_20_DFFSR_58 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_31_DFFSR_18 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_6_DFFPOSX1_23 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_11_DFFSR_226 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_6_OAI21X1_41 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_5_NAND2X1_59 DFFSR_62/gnd DFFSR_208/S FILL
XNAND2X1_56 INVX1_129/Y NAND2X1_57/B AND2X2_38/B NOR2X1_64/B DFFSR_59/S NAND2X1
XFILL_4_NAND2X1_62 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_5_OAI21X1_44 DFFSR_62/gnd DFFSR_208/S FILL
XOAI21X1_41 OAI21X1_41/A OAI21X1_41/B INVX1_152/A DFFSR_34/gnd OAI21X1_41/Y DFFSR_34/S
+ OAI21X1
XFILL_3_NAND2X1_65 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_3_DFFSR_113 BUFX2_99/A DFFSR_92/S FILL
XFILL_4_OAI21X1_47 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_0_OAI22X1_6 BUFX2_98/A DFFSR_32/S FILL
XFILL_44_DFFSR_144 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_2_NAND2X1_68 AND2X2_38/B DFFSR_23/S FILL
XFILL_3_OAI21X1_50 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_15_DFFPOSX1_42 INVX1_39/gnd DFFSR_34/S FILL
XFILL_7_DFFSR_220 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_4_NAND2X1_119 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_34_DFFSR_147 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_48_DFFSR_251 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_1_NAND2X1_71 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_2_OAI21X1_53 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_11_AOI22X1_19 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_24_DFFSR_150 AND2X2_38/B DFFSR_23/S FILL
XFILL_0_NAND2X1_74 AND2X2_38/B DFFSR_59/S FILL
XFILL_1_OAI21X1_56 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_39_DFFSR_25 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_28_DFFSR_65 BUFX2_79/A DFFSR_7/S FILL
XFILL_10_AOI22X1_22 INVX1_3/gnd DFFSR_79/S FILL
XFILL_0_INVX1_197 INVX1_3/gnd DFFSR_79/S FILL
XFILL_0_INVX1_59 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_38_DFFSR_254 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_14_DFFSR_153 INVX1_67/gnd DFFSR_201/S FILL
XFILL_0_OAI21X1_59 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_28_DFFSR_257 INVX1_39/gnd DFFSR_34/S FILL
XFILL_2_OAI21X1_101 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_18_DFFSR_260 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_25_DFFPOSX1_31 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_12_DFFSR_15 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_9_AOI22X1_25 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_8_AOI22X1_28 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_0_NAND3X1_179 NOR3X1_6/gnd DFFSR_79/S FILL
XNOR2X1_3 NOR2X1_3/A NOR2X1_3/B XOR2X1_4/gnd NOR2X1_3/Y DFFSR_91/S NOR2X1
XDFFSR_260 DFFSR_4/D CLKBUF1_4/Y DFFSR_257/R DFFSR_260/S DFFSR_260/D BUFX2_77/gnd
+ DFFSR_5/S DFFSR
XFILL_0_DFFSR_150 AND2X2_38/B DFFSR_23/S FILL
XFILL_25_0_2 AND2X2_38/B DFFSR_23/S FILL
XFILL_41_DFFSR_181 INVX1_3/gnd DFFSR_79/S FILL
XFILL_47_DFFSR_32 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_3_INVX1_124 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_36_DFFSR_72 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_4_DFFSR_257 INVX1_39/gnd DFFSR_34/S FILL
XFILL_31_DFFSR_184 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_1_NAND3X1_113 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_6_NAND2X1_20 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_21_DFFSR_187 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_3_DFFSR_29 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_20_DFFSR_22 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_3_NAND2X1_149 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_5_1_2 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_5_NAND2X1_23 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_11_DFFSR_190 INVX1_39/gnd DFFSR_34/S FILL
XNAND2X1_20 DFFSR_45/D AND2X2_5/Y DFFSR_8/gnd NAND3X1_36/A DFFSR_8/S NAND2X1
XFILL_4_NAND2X1_26 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_6_NOR2X1_66 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_3_NAND2X1_29 INVX1_3/gnd DFFSR_23/S FILL
XFILL_4_OAI21X1_11 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_9_DFFSR_4 DFFSR_4/gnd DFFSR_4/S FILL
XDFFPOSX1_23 NAND2X1_160/A CLKBUF1_45/Y AOI21X1_56/Y NOR3X1_6/gnd DFFSR_91/S DFFPOSX1
XFILL_44_DFFSR_108 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_2_NAND2X1_32 INVX1_3/gnd DFFSR_79/S FILL
XFILL_44_DFFSR_79 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_3_OAI21X1_14 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_7_DFFSR_184 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_34_DFFSR_111 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_5_10 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_9_NAND3X1_88 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_1_NAND2X1_35 INVX1_67/gnd DFFSR_201/S FILL
XFILL_48_DFFSR_215 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_2_OAI21X1_17 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_24_DFFSR_114 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_8_NAND3X1_91 AND2X2_38/B DFFSR_59/S FILL
XFILL_52_3_0 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_1_OAI21X1_20 AND2X2_38/B DFFSR_23/S FILL
XFILL_0_NAND2X1_38 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_28_DFFSR_29 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_38_DFFSR_218 BUFX2_98/A DFFSR_32/S FILL
XFILL_0_DFFSR_76 BUFX2_79/A DFFSR_7/S FILL
XFILL_0_INVX1_23 BUFX2_99/A DFFSR_7/S FILL
XFILL_0_INVX1_161 INVX1_1/gnd DFFSR_53/S FILL
XFILL_17_DFFSR_69 BUFX2_98/A DFFSR_32/S FILL
XFILL_3_AND2X2_28 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_14_DFFSR_117 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_7_NAND3X1_94 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_0_OAI21X1_23 INVX1_67/gnd DFFSR_201/S FILL
XFILL_28_DFFSR_221 AND2X2_38/B DFFSR_59/S FILL
XFILL_7_OR2X2_4 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_6_NAND3X1_97 AND2X2_38/B DFFSR_59/S FILL
XFILL_18_DFFSR_224 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_50_5_1 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_4_XOR2X1_6 BUFX2_99/A DFFSR_7/S FILL
XFILL_0_NAND3X1_143 BUFX2_8/gnd DFFSR_51/S FILL
XNAND3X1_97 DFFSR_173/Q BUFX2_30/Y BUFX2_26/Y AND2X2_38/B NAND3X1_97/Y DFFSR_59/S
+ NAND3X1
XFILL_9_NAND3X1_198 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_33_DFFSR_8 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_7_OAI22X1_4 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_5_DFFPOSX1_17 BUFX2_8/gnd DFFSR_51/S FILL
XDFFSR_224 DFFSR_224/Q CLKBUF1_10/Y BUFX2_64/Y DFFSR_151/S DFFSR_216/Q BUFX2_7/gnd
+ DFFSR_151/S DFFSR
XFILL_0_DFFSR_114 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_2_NAND2X1_179 INVX1_1/gnd DFFSR_97/S FILL
XFILL_41_DFFSR_145 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_30_1 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_8_DFFSR_83 INVX1_3/gnd DFFSR_79/S FILL
XFILL_36_DFFSR_36 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_25_DFFSR_76 BUFX2_79/A DFFSR_7/S FILL
XFILL_4_DFFSR_221 AND2X2_38/B DFFSR_59/S FILL
XFILL_31_DFFSR_148 INVX1_67/gnd DFFSR_175/S FILL
XFILL_45_DFFSR_252 AND2X2_38/B DFFSR_23/S FILL
XFILL_21_DFFSR_151 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_14_DFFPOSX1_36 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_35_DFFSR_255 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_3_NAND2X1_113 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_11_DFFSR_154 BUFX2_99/A DFFSR_7/S FILL
XFILL_25_DFFSR_258 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_2_AOI22X1_10 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_6_NOR2X1_30 INVX1_3/gnd DFFSR_23/S FILL
XFILL_15_DFFSR_261 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_16_6_0 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_1_AOI22X1_13 AND2X2_38/B DFFSR_23/S FILL
XFILL_11_OAI22X1_31 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_0_AOI22X1_16 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_10_OAI22X1_34 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_44_DFFSR_43 BUFX2_98/A DFFSR_6/S FILL
XFILL_33_DFFSR_83 INVX1_3/gnd DFFSR_79/S FILL
XFILL_7_DFFSR_148 INVX1_67/gnd DFFSR_175/S FILL
XFILL_24_DFFPOSX1_25 BUFX2_79/A DFFSR_6/S FILL
XFILL_48_DFFSR_179 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_8_NAND3X1_55 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_9_OAI22X1_37 INVX1_3/gnd DFFSR_23/S FILL
XFILL_0_DFFSR_40 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_8_NAND3X1_228 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_0_INVX1_125 AND2X2_38/B DFFSR_59/S FILL
XFILL_38_DFFSR_182 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_17_DFFSR_33 BUFX2_98/A DFFSR_32/S FILL
XFILL_7_NAND3X1_58 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_1_DFFSR_258 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_8_OAI22X1_40 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_4_BUFX2_68 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_4_DFFPOSX1_47 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_28_DFFSR_185 INVX1_39/gnd DFFSR_54/S FILL
XFILL_6_NAND3X1_61 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_7_OAI22X1_43 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_18_DFFSR_188 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_5_NAND3X1_64 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_6_OAI22X1_46 OR2X2_1/gnd DFFSR_59/S FILL
XNAND3X1_61 DFFSR_16/Q BUFX2_19/Y BUFX2_14/Y DFFSR_28/gnd NAND3X1_61/Y DFFSR_3/S NAND3X1
XFILL_0_NAND3X1_107 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_10_XOR2X1_3 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_4_NAND3X1_67 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_5_OAI22X1_49 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_41_DFFSR_90 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_3_NOR2X1_67 INVX1_67/gnd DFFSR_175/S FILL
XOAI22X1_46 INVX1_111/Y OAI22X1_43/B INVX1_112/Y OAI22X1_43/D OR2X2_1/gnd NOR2X1_56/B
+ DFFSR_59/S OAI22X1
XFILL_3_NAND3X1_70 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_4_OAI22X1_52 DFFSR_28/gnd DFFSR_3/S FILL
XDFFSR_188 INVX1_84/A DFFSR_1/CLK BUFX2_68/Y DFFSR_54/S DFFSR_172/Q DFFSR_46/gnd DFFSR_54/S
+ DFFSR
XFILL_2_NAND2X1_143 INVX1_67/gnd DFFSR_201/S FILL
XFILL_41_DFFSR_109 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_8_DFFSR_47 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_2_NAND3X1_73 INVX1_1/gnd DFFSR_97/S FILL
XFILL_25_DFFSR_40 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_14_DFFSR_80 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_4_DFFSR_185 INVX1_39/gnd DFFSR_54/S FILL
XFILL_31_DFFSR_112 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_1_NAND3X1_76 INVX1_1/gnd DFFSR_53/S FILL
XFILL_45_DFFSR_216 BUFX2_7/gnd DFFSR_216/S FILL
XNAND2X1_9 DFFSR_105/Q NOR2X1_5/Y BUFX2_79/A OAI21X1_1/C DFFSR_6/S NAND2X1
XFILL_21_DFFSR_115 INVX1_1/gnd DFFSR_97/S FILL
XFILL_0_NAND3X1_79 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_35_DFFSR_219 INVX1_67/gnd DFFSR_175/S FILL
XFILL_0_AND2X2_29 AND2X2_38/B DFFSR_23/S FILL
XFILL_11_DFFSR_118 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_26_1_0 INVX1_3/gnd DFFSR_23/S FILL
XFILL_4_NAND2X1_6 BUFX2_98/A DFFSR_32/S FILL
XFILL_25_DFFSR_222 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_49_DFFSR_97 INVX1_1/gnd DFFSR_97/S FILL
XFILL_15_DFFSR_225 INVX1_67/gnd DFFSR_175/S FILL
XFILL_20_DFFSR_2 BUFX2_79/A DFFSR_7/S FILL
XFILL_24_3_1 AND2X2_38/B DFFSR_59/S FILL
XOAI22X1_8 INVX1_19/Y OAI22X1_2/B INVX1_20/Y OAI22X1_2/D NOR3X1_6/gnd OAI22X1_8/Y
+ DFFSR_91/S OAI22X1
XINVX1_81 INVX1_81/A OR2X2_1/gnd INVX1_81/Y DFFSR_51/S INVX1
XFILL_33_DFFSR_47 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_5_DFFSR_94 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_22_DFFSR_87 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_7_DFFSR_112 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_6_2_0 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_4_OAI22X1_5 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_48_DFFSR_143 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_22_5_2 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_8_NAND3X1_19 BUFX2_99/A DFFSR_92/S FILL
XFILL_4_BUFX2_3 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_38_DFFSR_146 BUFX2_79/A DFFSR_7/S FILL
XFILL_8_NAND3X1_192 OR2X2_2/gnd DFFSR_216/S FILL
XINVX1_199 BUFX2_71/A DFFSR_62/gnd INVX1_199/Y DFFSR_62/S INVX1
XFILL_1_DFFSR_222 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_4_4_1 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_7_NAND3X1_22 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_4_BUFX2_32 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_28_DFFSR_149 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_4_DFFPOSX1_11 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_1_NAND2X1_173 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_6_NAND3X1_25 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_42_DFFSR_253 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_52_1 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_18_DFFSR_152 INVX1_1/gnd DFFSR_53/S FILL
XFILL_32_DFFSR_256 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_2_6_2 INVX1_67/gnd DFFSR_201/S FILL
XFILL_5_NAND3X1_28 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_6_OAI22X1_10 DFFSR_8/gnd DFFSR_60/S FILL
XNAND3X1_25 DFFSR_60/D BUFX2_17/Y BUFX2_12/Y DFFSR_8/gnd NAND3X1_25/Y DFFSR_8/S NAND3X1
XFILL_22_DFFSR_259 BUFX2_79/A DFFSR_6/S FILL
XFILL_4_NAND3X1_31 BUFX2_79/A DFFSR_6/S FILL
XFILL_5_OAI22X1_13 INVX1_1/gnd DFFSR_53/S FILL
XFILL_9_NAND3X1_126 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_2_INVX1_88 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_30_DFFSR_94 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_41_DFFSR_54 INVX1_39/gnd DFFSR_54/S FILL
XFILL_3_NOR2X1_31 INVX1_39/gnd DFFSR_54/S FILL
XOAI22X1_10 INVX1_24/Y OAI22X1_7/B INVX1_25/Y OAI22X1_7/D DFFSR_8/gnd NOR2X1_15/B
+ DFFSR_60/S OAI22X1
XFILL_13_DFFPOSX1_30 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_12_DFFSR_262 BUFX2_98/A DFFSR_32/S FILL
XFILL_3_NAND3X1_34 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_4_OAI22X1_16 AND2X2_38/B DFFSR_59/S FILL
XDFFSR_152 INVX1_115/A CLKBUF1_39/Y BUFX2_63/Y DFFSR_53/S DFFSR_160/Q INVX1_1/gnd
+ DFFSR_53/S DFFSR
XFILL_2_NAND2X1_107 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_3_OAI22X1_19 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_2_NAND3X1_37 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_8_DFFSR_11 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_14_DFFSR_44 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_4_DFFSR_149 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_1_BUFX2_79 BUFX2_79/A DFFSR_7/S FILL
XFILL_2_OAI22X1_22 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_1_NAND3X1_40 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_45_DFFSR_180 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_8_DFFSR_256 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_0_NAND3X1_43 BUFX2_99/A DFFSR_7/S FILL
XFILL_1_OAI22X1_25 INVX1_39/gnd DFFSR_54/S FILL
XFILL_35_DFFSR_183 INVX1_67/gnd DFFSR_175/S FILL
XFILL_23_DFFPOSX1_19 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_0_OAI22X1_28 INVX1_3/gnd DFFSR_23/S FILL
XFILL_25_DFFSR_186 BUFX2_99/A DFFSR_92/S FILL
XFILL_49_DFFSR_61 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_15_DFFSR_189 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_7_NAND3X1_222 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_3_DFFPOSX1_41 DFFSR_8/gnd DFFSR_60/S FILL
XINVX1_45 DFFSR_15/D OR2X2_3/gnd INVX1_45/Y DFFSR_4/S INVX1
XDFFSR_98 DFFSR_98/Q DFFSR_82/CLK DFFSR_5/R DFFSR_98/S DFFSR_98/D BUFX2_77/gnd DFFSR_98/S
+ DFFSR
XFILL_32_0_2 INVX1_1/gnd DFFSR_97/S FILL
XFILL_5_DFFSR_58 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_33_DFFSR_11 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_11_DFFSR_91 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_22_DFFSR_51 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_0_NOR2X1_68 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_48_DFFSR_107 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_38_DFFSR_110 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_8_NAND3X1_156 OR2X2_1/gnd DFFSR_59/S FILL
XINVX1_163 INVX1_163/A INVX1_39/gnd INVX1_163/Y DFFSR_54/S INVX1
XFILL_1_DFFSR_186 BUFX2_99/A DFFSR_92/S FILL
XFILL_28_DFFSR_113 BUFX2_99/A DFFSR_92/S FILL
XFILL_1_NAND2X1_137 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_42_DFFSR_217 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_4_INVX1_160 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_7_AND2X2_27 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_18_DFFSR_116 INVX1_3/gnd DFFSR_23/S FILL
XFILL_32_DFFSR_220 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_1_NAND2X1_7 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_22_DFFSR_223 INVX1_39/gnd DFFSR_34/S FILL
XFILL_30_DFFSR_58 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_2_INVX1_52 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_19_DFFSR_98 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_41_DFFSR_18 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_12_DFFSR_226 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_22_DFFPOSX1_49 BUFX2_99/A DFFSR_92/S FILL
XDFFSR_116 INVX1_30/A CLKBUF1_8/Y DFFSR_7/R DFFSR_23/S DFFSR_116/D INVX1_3/gnd DFFSR_23/S
+ DFFSR
XFILL_4_DFFSR_113 BUFX2_99/A DFFSR_92/S FILL
XFILL_1_BUFX2_43 AND2X2_38/B DFFSR_23/S FILL
XFILL_1_OAI22X1_6 BUFX2_98/A DFFSR_32/S FILL
XFILL_45_DFFSR_144 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_8_DFFSR_220 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_8_DFFSR_1 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_35_DFFSR_147 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_49_DFFSR_251 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_11_DFFSR_9 BUFX2_79/A DFFSR_6/S FILL
XFILL_25_DFFSR_150 AND2X2_38/B DFFSR_23/S FILL
XFILL_49_DFFSR_25 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_1_INVX1_197 INVX1_3/gnd DFFSR_79/S FILL
XFILL_39_DFFSR_254 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_38_DFFSR_65 BUFX2_79/A DFFSR_7/S FILL
XFILL_15_DFFSR_153 INVX1_67/gnd DFFSR_201/S FILL
XFILL_7_NAND3X1_186 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_29_DFFSR_257 INVX1_39/gnd DFFSR_34/S FILL
XFILL_19_DFFSR_260 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_0_NAND2X1_167 OR2X2_1/gnd DFFSR_59/S FILL
XDFFSR_62 DFFSR_62/Q CLKBUF1_31/Y DFFSR_1/R DFFSR_62/S DFFSR_62/D DFFSR_62/gnd DFFSR_62/S
+ DFFSR
XFILL_5_DFFSR_22 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_22_DFFSR_15 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_11_DFFSR_55 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_0_NOR2X1_32 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_6_OR2X2_1 OR2X2_1/gnd DFFSR_59/S FILL
XINVX1_127 NOR3X1_3/A BUFX2_8/gnd INVX1_127/Y DFFSR_51/S INVX1
XFILL_8_NAND3X1_120 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_4_NOR2X1_3 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_1_DFFSR_150 AND2X2_38/B DFFSR_23/S FILL
XFILL_12_DFFPOSX1_24 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_32_DFFSR_5 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_1_NAND2X1_101 INVX1_39/gnd DFFSR_54/S FILL
XFILL_42_DFFSR_181 INVX1_3/gnd DFFSR_79/S FILL
XFILL_46_DFFSR_72 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_5_DFFSR_257 INVX1_39/gnd DFFSR_34/S FILL
XFILL_32_DFFSR_184 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_23_6_0 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_22_DFFSR_187 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_30_DFFSR_22 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_2_DFFSR_69 BUFX2_98/A DFFSR_32/S FILL
XFILL_2_INVX1_16 BUFX2_99/A DFFSR_7/S FILL
XFILL_19_DFFSR_62 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_12_DFFSR_190 INVX1_39/gnd DFFSR_34/S FILL
XFILL_6_BUFX2_97 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_22_DFFPOSX1_13 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_6_NAND3X1_216 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_45_DFFSR_108 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_2_DFFPOSX1_35 INVX1_39/gnd DFFSR_54/S FILL
XFILL_8_DFFSR_184 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_35_DFFSR_111 DFFSR_8/gnd DFFSR_8/S FILL
XAND2X2_31 INVX1_135/A INVX1_145/A NOR3X1_6/gnd AND2X2_31/Y DFFSR_79/S AND2X2
XFILL_49_DFFSR_215 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_25_DFFSR_114 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_38_DFFSR_29 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_39_DFFSR_218 BUFX2_98/A DFFSR_32/S FILL
XFILL_1_INVX1_161 INVX1_1/gnd DFFSR_53/S FILL
XFILL_27_DFFSR_69 BUFX2_98/A DFFSR_32/S FILL
XFILL_4_AND2X2_28 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_15_DFFSR_117 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_7_NAND3X1_150 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_29_DFFSR_221 AND2X2_38/B DFFSR_59/S FILL
XFILL_19_DFFSR_224 BUFX2_7/gnd DFFSR_151/S FILL
XDFFSR_26 DFFSR_18/D DFFSR_92/CLK DFFSR_2/R DFFSR_6/S DFFSR_2/Q BUFX2_79/A DFFSR_6/S
+ DFFSR
XFILL_0_NAND2X1_131 INVX1_3/gnd DFFSR_79/S FILL
XFILL_11_DFFSR_19 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_8_OAI22X1_4 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_1_DFFSR_114 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_17_3 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_21_DFFPOSX1_43 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_33_1_0 INVX1_1/gnd DFFSR_53/S FILL
XFILL_42_DFFSR_145 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_46_DFFSR_36 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_35_DFFSR_76 BUFX2_79/A DFFSR_7/S FILL
XFILL_5_DFFSR_221 AND2X2_38/B DFFSR_59/S FILL
XFILL_32_DFFSR_148 INVX1_67/gnd DFFSR_175/S FILL
XFILL_5_NAND3X1_246 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_46_DFFSR_252 AND2X2_38/B DFFSR_23/S FILL
XFILL_22_DFFSR_151 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_31_3_1 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_36_DFFSR_255 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_2_DFFSR_33 BUFX2_98/A DFFSR_32/S FILL
XFILL_19_DFFSR_26 BUFX2_79/A DFFSR_6/S FILL
XFILL_12_DFFSR_154 BUFX2_99/A DFFSR_7/S FILL
XFILL_6_BUFX2_61 AND2X2_38/B DFFSR_59/S FILL
XFILL_26_DFFSR_258 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_8_OAI21X1_102 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_29_5_2 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_16_DFFSR_261 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_20_CLKBUF1_16 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_6_NAND3X1_180 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_19_CLKBUF1_19 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_8_DFFSR_148 INVX1_67/gnd DFFSR_175/S FILL
XFILL_43_DFFSR_83 INVX1_3/gnd DFFSR_79/S FILL
XFILL_18_CLKBUF1_22 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_49_DFFSR_179 OR2X2_1/gnd DFFSR_51/S FILL
XNAND3X1_216 NAND3X1_187/Y NAND3X1_219/B NAND3X1_215/Y DFFSR_46/gnd NAND3X1_216/Y
+ DFFSR_62/S NAND3X1
XFILL_9_6_2 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_17_CLKBUF1_25 INVX1_67/gnd DFFSR_201/S FILL
XFILL_1_INVX1_125 AND2X2_38/B DFFSR_59/S FILL
XFILL_39_DFFSR_182 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_27_DFFSR_33 BUFX2_98/A DFFSR_32/S FILL
XFILL_16_DFFSR_73 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_7_NAND3X1_114 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_2_DFFSR_258 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_16_CLKBUF1_28 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_29_DFFSR_185 INVX1_39/gnd DFFSR_54/S FILL
XFILL_11_DFFPOSX1_18 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_15_CLKBUF1_31 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_19_DFFSR_188 DFFSR_46/gnd DFFSR_54/S FILL
XNOR2X1_70 NOR2X1_70/A NOR2X1_70/B XOR2X1_4/gnd NOR2X1_70/Y DFFSR_91/S NOR2X1
XFILL_14_CLKBUF1_34 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_4_NOR2X1_67 INVX1_67/gnd DFFSR_175/S FILL
XFILL_13_CLKBUF1_37 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_12_CLKBUF1_40 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_42_DFFSR_109 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_35_DFFSR_40 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_24_DFFSR_80 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_7_DFFSR_87 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_11_CLKBUF1_43 AND2X2_38/B DFFSR_23/S FILL
XFILL_5_DFFSR_185 INVX1_39/gnd DFFSR_54/S FILL
XFILL_32_DFFSR_112 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_46_DFFSR_216 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_10_CLKBUF1_46 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_5_NAND3X1_210 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_22_DFFSR_115 INVX1_1/gnd DFFSR_97/S FILL
XFILL_1_DFFPOSX1_29 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_36_DFFSR_219 INVX1_67/gnd DFFSR_175/S FILL
XFILL_39_0_2 BUFX2_79/A DFFSR_6/S FILL
XFILL_1_AND2X2_29 AND2X2_38/B DFFSR_23/S FILL
XFILL_12_DFFSR_118 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_6_BUFX2_25 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_5_NAND2X1_6 BUFX2_98/A DFFSR_32/S FILL
XFILL_26_DFFSR_222 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_9_CLKBUF1_49 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_16_DFFSR_225 INVX1_67/gnd DFFSR_175/S FILL
XFILL_44_DFFSR_8 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_16_NOR3X1_4 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_6_NAND3X1_144 AND2X2_38/B DFFSR_59/S FILL
XFILL_10_DFFPOSX1_48 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_32_DFFSR_87 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_43_DFFSR_47 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_8_DFFSR_112 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_5_OAI22X1_5 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_49_DFFSR_143 OR2X2_2/gnd DFFSR_216/S FILL
XNAND3X1_180 AOI21X1_28/C AOI21X1_27/B AOI21X1_27/A OR2X2_1/gnd AOI21X1_21/B DFFSR_59/S
+ NAND3X1
XFILL_39_DFFSR_146 BUFX2_79/A DFFSR_7/S FILL
XFILL_16_DFFSR_37 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_2_DFFSR_222 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_3_BUFX2_72 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_29_DFFSR_149 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_39_3 BUFX2_79/A DFFSR_7/S FILL
XFILL_43_DFFSR_253 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_20_DFFPOSX1_37 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_19_DFFSR_152 INVX1_1/gnd DFFSR_53/S FILL
XFILL_33_DFFSR_256 DFFSR_8/gnd DFFSR_60/S FILL
XNOR2X1_34 NOR3X1_4/C NOR2X1_34/B XOR2X1_4/gnd NOR2X1_34/Y DFFSR_91/S NOR2X1
XFILL_23_DFFSR_259 BUFX2_79/A DFFSR_6/S FILL
XFILL_4_NAND3X1_240 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_40_DFFSR_94 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_51_DFFSR_54 INVX1_39/gnd DFFSR_54/S FILL
XFILL_4_NOR2X1_31 INVX1_39/gnd DFFSR_54/S FILL
XFILL_13_DFFSR_262 BUFX2_98/A DFFSR_32/S FILL
XFILL_1_AND2X2_3 INVX1_1/gnd DFFSR_53/S FILL
XFILL_24_DFFSR_44 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_7_DFFSR_51 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_5_DFFSR_149 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_13_DFFSR_84 BUFX2_99/A DFFSR_7/S FILL
XFILL_10_CLKBUF1_10 INVX1_67/gnd DFFSR_201/S FILL
XFILL_5_NAND3X1_174 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_46_DFFSR_180 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_9_DFFSR_256 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_36_DFFSR_183 INVX1_67/gnd DFFSR_175/S FILL
XFILL_26_DFFSR_186 BUFX2_99/A DFFSR_92/S FILL
XFILL_9_CLKBUF1_13 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_10_DFFSR_6 BUFX2_79/A DFFSR_6/S FILL
XFILL_16_DFFSR_189 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_8_CLKBUF1_16 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_6_NAND3X1_108 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_7_CLKBUF1_19 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_10_DFFPOSX1_12 AND2X2_38/B DFFSR_23/S FILL
XFILL_4_DFFSR_98 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_21_DFFSR_91 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_32_DFFSR_51 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_43_DFFSR_11 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_1_NOR2X1_68 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_6_CLKBUF1_22 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_49_DFFSR_107 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_5_CLKBUF1_25 INVX1_67/gnd DFFSR_201/S FILL
XNAND3X1_144 INVX1_144/A OAI21X1_32/Y OAI21X1_33/Y AND2X2_38/B AOI21X1_12/A DFFSR_59/S
+ NAND3X1
XFILL_30_6_0 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_39_DFFSR_110 OR2X2_3/gnd DFFSR_4/S FILL
XCLKBUF1_22 BUFX2_6/Y OR2X2_1/gnd CLKBUF1_22/Y DFFSR_59/S CLKBUF1
XOR2X2_2 OR2X2_2/A OR2X2_2/B OR2X2_2/gnd OR2X2_2/Y DFFSR_216/S OR2X2
XFILL_4_CLKBUF1_28 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_2_DFFSR_186 BUFX2_99/A DFFSR_92/S FILL
XFILL_3_BUFX2_36 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_29_DFFSR_113 BUFX2_99/A DFFSR_92/S FILL
XFILL_43_DFFSR_217 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_3_CLKBUF1_31 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_8_AND2X2_27 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_19_DFFSR_116 INVX1_3/gnd DFFSR_23/S FILL
XFILL_2_CLKBUF1_34 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_33_DFFSR_220 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_31_DFFSR_2 BUFX2_79/A DFFSR_7/S FILL
XFILL_2_NAND2X1_7 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_23_DFFSR_223 INVX1_39/gnd DFFSR_34/S FILL
XFILL_1_CLKBUF1_37 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_4_NAND3X1_204 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_40_DFFSR_58 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_1_INVX1_92 AND2X2_38/B DFFSR_23/S FILL
XFILL_29_DFFSR_98 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_13_DFFSR_226 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_0_CLKBUF1_40 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_0_DFFPOSX1_23 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_7_DFFSR_15 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_13_DFFSR_48 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_5_DFFSR_113 BUFX2_99/A DFFSR_92/S FILL
XFILL_2_OAI22X1_6 BUFX2_98/A DFFSR_32/S FILL
XFILL_0_BUFX2_83 BUFX2_79/A DFFSR_7/S FILL
XFILL_5_NAND3X1_138 INVX1_67/gnd DFFSR_201/S FILL
XFILL_46_DFFSR_144 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_9_DFFSR_220 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_36_DFFSR_147 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_50_DFFSR_251 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_26_DFFSR_150 AND2X2_38/B DFFSR_23/S FILL
XFILL_2_INVX1_197 INVX1_3/gnd DFFSR_79/S FILL
XFILL_40_DFFSR_254 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_48_DFFSR_65 BUFX2_79/A DFFSR_7/S FILL
XFILL_16_DFFSR_153 INVX1_67/gnd DFFSR_201/S FILL
XFILL_30_DFFSR_257 INVX1_39/gnd DFFSR_34/S FILL
XFILL_20_DFFSR_260 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_32_DFFSR_15 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_21_DFFSR_55 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_10_DFFSR_95 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_40_1_0 BUFX2_98/A DFFSR_6/S FILL
XFILL_19_DFFPOSX1_31 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_4_DFFSR_62 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_1_NOR2X1_32 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_10_DFFSR_263 OR2X2_1/gnd DFFSR_51/S FILL
XNAND3X1_108 NAND2X1_48/Y NAND3X1_105/Y AND2X2_24/Y BUFX2_8/gnd NOR2X1_52/A DFFSR_81/S
+ NAND3X1
XFILL_3_NAND3X1_234 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_38_3_1 BUFX2_79/A DFFSR_7/S FILL
XFILL_2_DFFSR_150 AND2X2_38/B DFFSR_23/S FILL
XFILL_43_DFFSR_181 INVX1_3/gnd DFFSR_79/S FILL
XFILL_6_DFFSR_257 INVX1_39/gnd DFFSR_34/S FILL
XFILL_33_DFFSR_184 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_36_5_2 BUFX2_99/A DFFSR_92/S FILL
XFILL_23_DFFSR_187 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_4_NAND3X1_168 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_40_DFFSR_22 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_1_INVX1_56 BUFX2_98/A DFFSR_6/S FILL
XFILL_29_DFFSR_62 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_13_DFFSR_190 INVX1_39/gnd DFFSR_34/S FILL
XFILL_9_DFFPOSX1_42 INVX1_39/gnd DFFSR_34/S FILL
XFILL_13_DFFSR_12 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_0_BUFX2_47 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_46_DFFSR_108 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_5_NAND3X1_102 INVX1_3/gnd DFFSR_23/S FILL
XFILL_9_DFFSR_184 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_36_DFFSR_111 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_50_DFFSR_215 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_26_DFFSR_114 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_40_DFFSR_218 BUFX2_98/A DFFSR_32/S FILL
XFILL_2_INVX1_161 INVX1_1/gnd DFFSR_53/S FILL
XFILL_48_DFFSR_29 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_37_DFFSR_69 BUFX2_98/A DFFSR_32/S FILL
XFILL_5_AND2X2_28 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_16_DFFSR_117 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_30_DFFSR_221 AND2X2_38/B DFFSR_59/S FILL
XFILL_20_DFFSR_224 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_4_DFFSR_26 BUFX2_79/A DFFSR_6/S FILL
XFILL_21_DFFSR_19 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_10_DFFSR_59 AND2X2_38/B DFFSR_59/S FILL
XFILL_10_DFFSR_227 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_3_NAND3X1_198 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_9_OAI22X1_4 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_3_NOR2X1_7 BUFX2_98/A DFFSR_32/S FILL
XFILL_2_DFFSR_114 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_46_0_2 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_22_DFFSR_9 BUFX2_79/A DFFSR_6/S FILL
XFILL_43_DFFSR_145 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_45_DFFSR_76 BUFX2_79/A DFFSR_7/S FILL
XFILL_6_DFFSR_221 AND2X2_38/B DFFSR_59/S FILL
XFILL_33_DFFSR_148 INVX1_67/gnd DFFSR_175/S FILL
XFILL_47_DFFSR_252 AND2X2_38/B DFFSR_23/S FILL
XFILL_23_DFFSR_151 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_4_NAND3X1_132 AND2X2_38/B DFFSR_23/S FILL
XFILL_37_DFFSR_255 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_29_DFFSR_26 BUFX2_79/A DFFSR_6/S FILL
XFILL_1_INVX1_20 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_1_DFFSR_73 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_18_DFFSR_66 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_13_DFFSR_154 BUFX2_99/A DFFSR_7/S FILL
XFILL_27_DFFSR_258 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_6_NAND2X1_168 BUFX2_79/A DFFSR_6/S FILL
XFILL_17_DFFSR_261 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_0_BUFX2_11 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_5_XOR2X1_3 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_21_DFFPOSX1_1 INVX1_39/gnd DFFSR_34/S FILL
XFILL_9_DFFSR_148 INVX1_67/gnd DFFSR_175/S FILL
XFILL_43_DFFSR_5 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_20_DFFPOSX1_4 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_18_DFFPOSX1_25 BUFX2_79/A DFFSR_6/S FILL
XFILL_50_DFFSR_179 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_19_DFFPOSX1_7 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_12_1_1 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_2_INVX1_125 AND2X2_38/B DFFSR_59/S FILL
XFILL_40_DFFSR_182 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_9_DFFSR_80 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_37_DFFSR_33 BUFX2_98/A DFFSR_32/S FILL
XFILL_26_DFFSR_73 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_2_NAND3X1_228 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_3_DFFSR_258 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_30_DFFSR_185 INVX1_39/gnd DFFSR_54/S FILL
XFILL_20_DFFSR_188 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_10_3_2 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_10_DFFSR_23 AND2X2_38/B DFFSR_23/S FILL
XFILL_10_DFFSR_191 INVX1_67/gnd DFFSR_175/S FILL
XFILL_5_NOR2X1_67 INVX1_67/gnd DFFSR_175/S FILL
XFILL_3_NAND3X1_162 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_1_NOR3X1_4 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_8_DFFPOSX1_36 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_43_DFFSR_109 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_45_DFFSR_40 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_34_DFFSR_80 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_6_DFFSR_185 INVX1_39/gnd DFFSR_54/S FILL
XFILL_33_DFFSR_112 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_47_DFFSR_216 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_23_DFFSR_115 INVX1_1/gnd DFFSR_97/S FILL
XFILL_37_DFFSR_219 INVX1_67/gnd DFFSR_175/S FILL
XFILL_1_DFFSR_37 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_18_DFFSR_30 BUFX2_98/A DFFSR_32/S FILL
XFILL_2_AND2X2_29 AND2X2_38/B DFFSR_23/S FILL
XFILL_13_DFFSR_118 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_5_BUFX2_65 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_6_NAND2X1_6 BUFX2_98/A DFFSR_32/S FILL
XFILL_27_DFFSR_222 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_6_NAND2X1_132 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_17_DFFSR_225 INVX1_67/gnd DFFSR_175/S FILL
XFILL_37_6_0 BUFX2_99/A DFFSR_7/S FILL
XXOR2X1_7 XOR2X1_7/A XOR2X1_7/B BUFX2_98/A XOR2X1_7/Y DFFSR_6/S XOR2X1
XFILL_42_DFFSR_87 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_9_DFFSR_112 OR2X2_4/gnd DFFSR_32/S FILL
XNAND2X1_168 NAND2X1_167/B INVX1_208/Y BUFX2_79/A AOI21X1_60/A DFFSR_6/S NAND2X1
XFILL_6_OAI22X1_5 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_50_DFFSR_143 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_4_OAI21X1_114 AND2X2_38/B DFFSR_59/S FILL
XFILL_27_DFFPOSX1_44 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_8_AOI21X1_60 BUFX2_79/A DFFSR_7/S FILL
XFILL_40_DFFSR_146 BUFX2_79/A DFFSR_7/S FILL
XFILL_26_DFFSR_37 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_9_DFFSR_44 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_7_AOI21X1_63 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_2_NAND3X1_192 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_15_DFFSR_77 BUFX2_98/A DFFSR_32/S FILL
XFILL_3_DFFSR_222 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_30_DFFSR_149 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_6_AOI21X1_66 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_44_DFFSR_253 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_20_DFFSR_152 INVX1_1/gnd DFFSR_53/S FILL
XFILL_34_DFFSR_256 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_5_AOI21X1_69 INVX1_1/gnd DFFSR_97/S FILL
XAOI21X1_66 AND2X2_42/Y AOI21X1_66/B NOR2X1_80/Y NOR3X1_6/gnd AOI21X1_66/Y DFFSR_91/S
+ AOI21X1
XFILL_10_DFFSR_155 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_24_DFFSR_259 BUFX2_79/A DFFSR_6/S FILL
XFILL_50_DFFSR_94 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_5_NOR2X1_31 INVX1_39/gnd DFFSR_54/S FILL
XFILL_3_NAND3X1_126 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_14_DFFSR_262 BUFX2_98/A DFFSR_32/S FILL
XFILL_5_NAND2X1_162 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_6_DFFSR_91 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_6_DFFSR_149 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_34_DFFSR_44 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_23_DFFSR_84 BUFX2_99/A DFFSR_7/S FILL
XFILL_47_DFFSR_180 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_37_DFFSR_183 INVX1_67/gnd DFFSR_175/S FILL
XBUFX2_69 BUFX2_60/A DFFSR_1/gnd BUFX2_69/Y DFFSR_1/S BUFX2
XFILL_47_1_0 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_0_DFFSR_259 BUFX2_79/A DFFSR_6/S FILL
XFILL_5_BUFX2_29 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_27_DFFSR_186 BUFX2_99/A DFFSR_92/S FILL
XFILL_17_DFFPOSX1_19 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_17_DFFSR_189 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_1_NAND3X1_222 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_9_DFFPOSX1_1 INVX1_39/gnd DFFSR_34/S FILL
XFILL_45_3_1 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_31_DFFSR_91 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_42_DFFSR_51 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_3_INVX1_85 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_8_DFFPOSX1_4 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_2_NOR2X1_68 OR2X2_2/gnd DFFSR_175/S FILL
XNAND2X1_132 DFFSR_265/Q DFFSR_151/S XOR2X1_1/gnd NAND2X1_132/Y DFFSR_151/S NAND2X1
XFILL_50_DFFSR_107 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_7_DFFPOSX1_7 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_8_AOI21X1_24 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_43_5_2 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_40_DFFSR_110 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_15_DFFSR_41 BUFX2_98/A DFFSR_6/S FILL
XFILL_7_AOI21X1_27 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_2_NAND3X1_156 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_3_DFFSR_186 BUFX2_99/A DFFSR_92/S FILL
XFILL_2_BUFX2_76 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_30_DFFSR_113 BUFX2_99/A DFFSR_92/S FILL
XFILL_6_AOI21X1_30 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_44_DFFSR_217 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_7_DFFPOSX1_30 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_20_DFFSR_116 INVX1_3/gnd DFFSR_23/S FILL
XFILL_5_AOI21X1_33 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_34_DFFSR_220 BUFX2_7/gnd DFFSR_151/S FILL
XAOI21X1_30 INVX1_160/Y AOI21X1_30/B NOR2X1_70/Y XOR2X1_4/gnd AOI21X1_30/Y DFFSR_97/S
+ AOI21X1
XFILL_10_DFFSR_119 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_3_NAND2X1_7 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_4_AOI21X1_36 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_24_DFFSR_223 INVX1_39/gnd DFFSR_34/S FILL
XFILL_50_DFFSR_58 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_39_DFFSR_98 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_3_AOI21X1_39 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_14_DFFSR_226 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_16_DFFPOSX1_49 BUFX2_99/A DFFSR_92/S FILL
XFILL_2_AOI21X1_42 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_11_4_0 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_0_AND2X2_7 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_5_NAND2X1_126 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_6_DFFSR_55 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_23_DFFSR_48 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_12_DFFSR_88 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_6_DFFSR_113 BUFX2_99/A DFFSR_92/S FILL
XFILL_1_AOI21X1_45 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_3_OAI22X1_6 BUFX2_98/A DFFSR_32/S FILL
XFILL_47_DFFSR_144 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_0_AOI21X1_48 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_37_DFFSR_147 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_51_DFFSR_251 BUFX2_7/gnd DFFSR_151/S FILL
XBUFX2_33 BUFX2_34/A NOR3X1_6/gnd BUFX2_33/Y DFFSR_91/S BUFX2
XFILL_0_DFFSR_223 INVX1_39/gnd DFFSR_34/S FILL
XFILL_27_DFFSR_150 AND2X2_38/B DFFSR_23/S FILL
XFILL_3_OAI21X1_108 INVX1_1/gnd DFFSR_53/S FILL
XFILL_26_DFFPOSX1_38 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_41_DFFSR_254 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_3_INVX1_197 INVX1_3/gnd DFFSR_79/S FILL
XFILL_17_DFFSR_153 INVX1_67/gnd DFFSR_201/S FILL
XFILL_48_5 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_8_OAI21X1_72 INVX1_3/gnd DFFSR_23/S FILL
XFILL_31_DFFSR_257 INVX1_39/gnd DFFSR_34/S FILL
XFILL_1_NAND3X1_186 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_6_NAND2X1_93 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_7_OAI21X1_75 INVX1_39/gnd DFFSR_54/S FILL
XFILL_21_DFFSR_260 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_53_0_2 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_42_DFFSR_15 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_31_DFFSR_55 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_3_INVX1_49 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_20_DFFSR_95 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_2_NOR2X1_32 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_6_OAI21X1_78 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_5_NAND2X1_96 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_11_DFFSR_263 OR2X2_1/gnd DFFSR_51/S FILL
XNAND2X1_93 AND2X2_34/B INVX1_159/A XOR2X1_4/gnd XOR2X1_4/B DFFSR_91/S NAND2X1
XFILL_5_OAI21X1_81 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_4_NAND2X1_99 INVX1_39/gnd DFFSR_54/S FILL
XOAI21X1_78 INVX1_167/A INVX1_168/A OAI21X1_78/C OR2X2_6/gnd INVX1_177/A DFFSR_92/S
+ OAI21X1
XFILL_2_NAND3X1_120 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_4_OAI21X1_84 BUFX2_98/A DFFSR_6/S FILL
XFILL_3_DFFSR_150 AND2X2_38/B DFFSR_23/S FILL
XFILL_2_BUFX2_40 INVX1_1/gnd DFFSR_97/S FILL
XFILL_44_DFFSR_181 INVX1_3/gnd DFFSR_79/S FILL
XFILL_3_OAI21X1_87 BUFX2_79/A DFFSR_7/S FILL
XFILL_7_DFFSR_257 INVX1_39/gnd DFFSR_34/S FILL
XFILL_4_NAND2X1_156 AND2X2_38/B DFFSR_59/S FILL
XFILL_34_DFFSR_184 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_2_OAI21X1_90 BUFX2_98/A DFFSR_32/S FILL
XFILL_21_DFFSR_6 BUFX2_79/A DFFSR_6/S FILL
XFILL_24_DFFSR_187 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_1_OAI21X1_93 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_50_DFFSR_22 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_0_INVX1_96 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_39_DFFSR_62 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_14_DFFSR_190 INVX1_39/gnd DFFSR_34/S FILL
XFILL_0_OAI21X1_96 AND2X2_38/B DFFSR_59/S FILL
XFILL_16_DFFPOSX1_13 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_6_DFFSR_19 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_5_BUFX2_7 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_23_DFFSR_12 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_12_DFFSR_52 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_19_1_1 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_47_DFFSR_108 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_0_NAND3X1_216 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_1_0_0 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_0_AOI21X1_12 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_37_DFFSR_111 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_17_3_2 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_0_DFFSR_187 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_27_DFFSR_114 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_42_DFFSR_2 BUFX2_79/A DFFSR_7/S FILL
XFILL_41_DFFSR_218 BUFX2_98/A DFFSR_32/S FILL
XFILL_3_INVX1_161 INVX1_1/gnd DFFSR_53/S FILL
XFILL_9_OAI21X1_33 INVX1_3/gnd DFFSR_79/S FILL
XFILL_47_DFFSR_69 BUFX2_98/A DFFSR_32/S FILL
XFILL_6_AND2X2_28 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_17_DFFSR_117 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_31_DFFSR_221 AND2X2_38/B DFFSR_59/S FILL
XFILL_8_OAI21X1_36 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_1_NAND3X1_150 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_0_NAND2X1_8 INVX1_1/gnd DFFSR_53/S FILL
XFILL_6_NAND2X1_57 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_7_OAI21X1_39 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_21_DFFSR_224 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_31_DFFSR_19 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_3_INVX1_13 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_3_DFFSR_66 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_20_DFFSR_59 AND2X2_38/B DFFSR_59/S FILL
XFILL_6_DFFPOSX1_24 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_6_OAI21X1_42 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_5_NAND2X1_60 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_11_DFFSR_227 BUFX2_7/gnd DFFSR_151/S FILL
XNAND2X1_57 INVX1_3/A NAND2X1_57/B DFFSR_1/gnd AOI21X1_6/B DFFSR_1/S NAND2X1
XFILL_4_NAND2X1_63 AND2X2_38/B DFFSR_59/S FILL
XFILL_5_OAI21X1_45 DFFSR_62/gnd DFFSR_208/S FILL
XOAI21X1_42 NOR3X1_5/B NOR3X1_5/C NOR3X1_5/A BUFX2_7/gnd OAI21X1_42/Y DFFSR_151/S
+ OAI21X1
XFILL_3_DFFSR_114 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_4_OAI21X1_48 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_3_NAND2X1_66 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_0_OAI22X1_7 AND2X2_38/B DFFSR_59/S FILL
XFILL_44_DFFSR_145 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_15_DFFPOSX1_43 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_2_NAND2X1_69 INVX1_3/gnd DFFSR_23/S FILL
XFILL_3_OAI21X1_51 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_7_DFFSR_221 AND2X2_38/B DFFSR_59/S FILL
XFILL_34_DFFSR_148 INVX1_67/gnd DFFSR_175/S FILL
XFILL_4_NAND2X1_120 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_1_NAND2X1_72 AND2X2_38/B DFFSR_59/S FILL
XFILL_2_OAI21X1_54 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_48_DFFSR_252 AND2X2_38/B DFFSR_23/S FILL
XFILL_11_AOI22X1_20 INVX1_39/gnd DFFSR_34/S FILL
XFILL_44_6_0 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_24_DFFSR_151 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_38_DFFSR_255 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_0_NAND2X1_75 INVX1_3/gnd DFFSR_79/S FILL
XFILL_1_OAI21X1_57 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_28_DFFSR_66 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_39_DFFSR_26 BUFX2_79/A DFFSR_6/S FILL
XFILL_0_INVX1_198 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_10_AOI22X1_23 INVX1_39/gnd DFFSR_34/S FILL
XFILL_0_INVX1_60 INVX1_39/gnd DFFSR_34/S FILL
XFILL_14_DFFSR_154 BUFX2_99/A DFFSR_7/S FILL
XFILL_0_OAI21X1_60 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_28_DFFSR_258 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_2_OAI21X1_102 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_25_DFFPOSX1_32 INVX1_67/gnd DFFSR_201/S FILL
XFILL_18_DFFSR_261 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_12_DFFSR_16 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_9_AOI22X1_26 INVX1_1/gnd DFFSR_97/S FILL
XFILL_0_NAND3X1_180 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_8_AOI22X1_29 INVX1_1/gnd DFFSR_53/S FILL
XNOR2X1_4 INVX1_3/A NOR3X1_1/A INVX1_1/gnd NOR2X1_4/Y DFFSR_53/S NOR2X1
XFILL_51_DFFSR_179 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_0_DFFSR_151 XOR2X1_1/gnd DFFSR_151/S FILL
XDFFSR_261 DFFSR_5/D DFFSR_5/CLK DFFSR_257/R DFFSR_98/S DFFSR_261/D BUFX2_77/gnd DFFSR_98/S
+ DFFSR
XFILL_3_INVX1_125 AND2X2_38/B DFFSR_59/S FILL
XFILL_41_DFFSR_182 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_47_DFFSR_33 BUFX2_98/A DFFSR_32/S FILL
XFILL_36_DFFSR_73 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_4_DFFSR_258 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_31_DFFSR_185 INVX1_39/gnd DFFSR_54/S FILL
XFILL_1_NAND3X1_114 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_6_NAND2X1_21 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_21_DFFSR_188 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_3_DFFSR_30 BUFX2_98/A DFFSR_32/S FILL
XFILL_20_DFFSR_23 AND2X2_38/B DFFSR_23/S FILL
XFILL_5_NAND2X1_24 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_11_DFFSR_191 INVX1_67/gnd DFFSR_175/S FILL
XFILL_3_NAND2X1_150 DFFSR_1/gnd DFFSR_1/S FILL
XNAND2X1_21 DFFSR_118/D NOR2X1_5/Y DFFSR_28/gnd OAI21X1_6/C DFFSR_8/S NAND2X1
XFILL_4_NAND2X1_27 AND2X2_38/B DFFSR_23/S FILL
XFILL_6_NOR2X1_67 INVX1_67/gnd DFFSR_175/S FILL
XFILL_8_1 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_9_DFFSR_5 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_3_NAND2X1_30 AND2X2_38/B DFFSR_23/S FILL
XFILL_4_OAI21X1_12 OR2X2_1/gnd DFFSR_51/S FILL
XDFFPOSX1_24 NAND2X1_165/B CLKBUF1_48/Y AOI21X1_59/Y BUFX2_8/gnd DFFSR_51/S DFFPOSX1
XFILL_44_DFFSR_109 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_54_1_0 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_2_NAND2X1_33 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_3_OAI21X1_15 INVX1_3/gnd DFFSR_79/S FILL
XFILL_44_DFFSR_80 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_7_DFFSR_185 INVX1_39/gnd DFFSR_54/S FILL
XFILL_34_DFFSR_112 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_1_NAND2X1_36 INVX1_3/gnd DFFSR_79/S FILL
XFILL_2_OAI21X1_18 INVX1_39/gnd DFFSR_34/S FILL
XFILL_48_DFFSR_216 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_24_DFFSR_115 INVX1_1/gnd DFFSR_97/S FILL
XFILL_8_NAND3X1_92 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_38_DFFSR_219 INVX1_67/gnd DFFSR_175/S FILL
XFILL_52_3_1 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_0_NAND2X1_39 BUFX2_98/A DFFSR_6/S FILL
XFILL_1_OAI21X1_21 AND2X2_38/B DFFSR_59/S FILL
XFILL_17_DFFSR_70 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_0_INVX1_24 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_28_DFFSR_30 BUFX2_98/A DFFSR_32/S FILL
XFILL_0_DFFSR_77 BUFX2_98/A DFFSR_32/S FILL
XFILL_0_INVX1_162 INVX1_39/gnd DFFSR_34/S FILL
XFILL_3_AND2X2_29 AND2X2_38/B DFFSR_23/S FILL
XFILL_14_DFFSR_118 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_7_NAND3X1_95 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_28_DFFSR_222 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_0_OAI21X1_24 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_6_NAND3X1_98 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_7_OR2X2_5 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_18_DFFSR_225 INVX1_67/gnd DFFSR_175/S FILL
XFILL_50_5_2 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_0_NAND3X1_144 AND2X2_38/B DFFSR_59/S FILL
XFILL_4_XOR2X1_7 BUFX2_98/A DFFSR_6/S FILL
XNAND3X1_98 DFFSR_157/D AND2X2_18/B BUFX2_29/Y OR2X2_1/gnd AND2X2_23/B DFFSR_59/S
+ NAND3X1
XFILL_33_DFFSR_9 BUFX2_79/A DFFSR_6/S FILL
XFILL_7_OAI22X1_5 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_51_DFFSR_143 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_5_DFFPOSX1_18 DFFSR_46/gnd DFFSR_62/S FILL
XDFFSR_225 DFFSR_225/Q CLKBUF1_34/Y BUFX2_62/Y DFFSR_175/S DFFSR_217/Q INVX1_67/gnd
+ DFFSR_175/S DFFSR
XFILL_2_NAND2X1_180 INVX1_1/gnd DFFSR_97/S FILL
XFILL_0_DFFSR_115 INVX1_1/gnd DFFSR_97/S FILL
XFILL_41_DFFSR_146 BUFX2_79/A DFFSR_7/S FILL
XFILL_30_2 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_36_DFFSR_37 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_8_DFFSR_84 BUFX2_99/A DFFSR_7/S FILL
XFILL_25_DFFSR_77 BUFX2_98/A DFFSR_32/S FILL
XFILL_4_DFFSR_222 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_31_DFFSR_149 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_45_DFFSR_253 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_21_DFFSR_152 INVX1_1/gnd DFFSR_53/S FILL
XFILL_14_DFFPOSX1_37 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_35_DFFSR_256 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_18_4_0 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_3_NAND2X1_114 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_11_DFFSR_155 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_2_AOI22X1_11 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_25_DFFSR_259 BUFX2_79/A DFFSR_6/S FILL
XFILL_6_NOR2X1_31 INVX1_39/gnd DFFSR_54/S FILL
XFILL_15_DFFSR_262 BUFX2_98/A DFFSR_32/S FILL
XFILL_16_6_1 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_1_AOI22X1_14 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_17_NOR3X1_1 INVX1_3/gnd DFFSR_79/S FILL
XFILL_11_OAI22X1_32 INVX1_39/gnd DFFSR_54/S FILL
XFILL_0_AOI22X1_17 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_10_OAI22X1_35 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_44_DFFSR_44 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_33_DFFSR_84 BUFX2_99/A DFFSR_7/S FILL
XFILL_7_DFFSR_149 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_24_DFFPOSX1_26 AND2X2_38/B DFFSR_23/S FILL
XFILL_9_NAND3X1_53 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_48_DFFSR_180 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_8_NAND3X1_56 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_9_OAI22X1_38 AND2X2_38/B DFFSR_23/S FILL
XFILL_38_DFFSR_183 INVX1_67/gnd DFFSR_175/S FILL
XFILL_8_NAND3X1_229 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_0_DFFSR_41 BUFX2_98/A DFFSR_6/S FILL
XFILL_0_INVX1_126 INVX1_3/gnd DFFSR_23/S FILL
XFILL_17_DFFSR_34 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_7_NAND3X1_59 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_1_DFFSR_259 BUFX2_79/A DFFSR_6/S FILL
XFILL_4_BUFX2_69 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_8_OAI22X1_41 INVX1_39/gnd DFFSR_54/S FILL
XFILL_28_DFFSR_186 BUFX2_99/A DFFSR_92/S FILL
XFILL_4_DFFPOSX1_48 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_6_NAND3X1_62 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_7_OAI22X1_44 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_18_DFFSR_189 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_5_NAND3X1_65 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_6_OAI22X1_47 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_0_NAND3X1_108 BUFX2_8/gnd DFFSR_81/S FILL
XNAND3X1_62 DFFSR_72/Q BUFX2_15/Y NOR2X1_2/Y DFFSR_8/gnd NAND3X1_63/B DFFSR_60/S NAND3X1
XFILL_10_XOR2X1_4 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_4_NAND3X1_68 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_41_DFFSR_91 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_5_OAI22X1_50 INVX1_3/gnd DFFSR_23/S FILL
XFILL_3_NOR2X1_68 OR2X2_2/gnd DFFSR_175/S FILL
XOAI22X1_47 INVX1_113/Y OAI22X1_41/B INVX1_114/Y OAI22X1_41/D BUFX2_8/gnd NOR2X1_56/A
+ DFFSR_81/S OAI22X1
XFILL_3_NAND3X1_71 BUFX2_7/gnd DFFSR_216/S FILL
XDFFSR_189 INVX1_91/A CLKBUF1_12/Y BUFX2_70/Y DFFSR_51/S DFFSR_173/Q BUFX2_8/gnd DFFSR_51/S
+ DFFSR
XFILL_2_NAND2X1_144 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_41_DFFSR_110 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_2_NAND3X1_74 INVX1_1/gnd DFFSR_97/S FILL
XFILL_8_DFFSR_48 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_25_DFFSR_41 BUFX2_98/A DFFSR_6/S FILL
XFILL_14_DFFSR_81 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_4_DFFSR_186 BUFX2_99/A DFFSR_92/S FILL
XFILL_31_DFFSR_113 BUFX2_99/A DFFSR_92/S FILL
XFILL_1_NAND3X1_77 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_45_DFFSR_217 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_21_DFFSR_116 INVX1_3/gnd DFFSR_23/S FILL
XFILL_0_NAND3X1_80 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_35_DFFSR_220 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_0_AND2X2_30 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_11_DFFSR_119 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_4_NAND2X1_7 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_26_1_1 INVX1_3/gnd DFFSR_23/S FILL
XFILL_25_DFFSR_223 INVX1_39/gnd DFFSR_34/S FILL
XFILL_49_DFFSR_98 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_8_0_0 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_15_DFFSR_226 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_20_DFFSR_3 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_24_3_2 AND2X2_38/B DFFSR_59/S FILL
XOAI22X1_9 INVX1_21/Y OAI22X1_6/B INVX1_22/Y OAI22X1_6/D OR2X2_4/gnd NOR2X1_13/A DFFSR_3/S
+ OAI22X1
XINVX1_82 INVX1_82/A XOR2X1_1/gnd INVX1_82/Y DFFSR_151/S INVX1
XFILL_33_DFFSR_48 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_22_DFFSR_88 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_5_DFFSR_95 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_7_DFFSR_113 BUFX2_99/A DFFSR_92/S FILL
XFILL_6_2_1 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_4_OAI22X1_6 BUFX2_98/A DFFSR_32/S FILL
XFILL_48_DFFSR_144 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_8_NAND3X1_20 BUFX2_99/A DFFSR_7/S FILL
XFILL_4_BUFX2_4 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_38_DFFSR_147 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_8_NAND3X1_193 XOR2X1_1/gnd DFFSR_208/S FILL
XINVX1_200 BUFX2_72/A BUFX2_72/gnd INVX1_200/Y DFFSR_201/S INVX1
XFILL_4_4_2 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_7_NAND3X1_23 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_4_BUFX2_33 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_1_DFFSR_223 INVX1_39/gnd DFFSR_34/S FILL
XFILL_28_DFFSR_150 AND2X2_38/B DFFSR_23/S FILL
XFILL_4_DFFPOSX1_12 AND2X2_38/B DFFSR_23/S FILL
XFILL_1_NAND2X1_174 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_42_DFFSR_254 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_6_NAND3X1_26 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_52_2 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_18_DFFSR_153 INVX1_67/gnd DFFSR_201/S FILL
XFILL_5_NAND3X1_29 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_32_DFFSR_257 INVX1_39/gnd DFFSR_34/S FILL
XFILL_6_OAI22X1_11 BUFX2_99/A DFFSR_92/S FILL
XNAND3X1_26 DFFSR_4/Q NOR2X1_4/Y BUFX2_17/Y DFFSR_28/gnd AND2X2_9/B DFFSR_3/S NAND3X1
XFILL_22_DFFSR_260 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_5_OAI22X1_14 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_41_DFFSR_55 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_4_NAND3X1_32 BUFX2_79/A DFFSR_7/S FILL
XFILL_2_INVX1_89 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_9_NAND3X1_127 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_30_DFFSR_95 DFFSR_5/gnd DFFSR_5/S FILL
XOAI22X1_11 INVX1_26/Y OAI22X1_2/B INVX1_27/Y OAI22X1_2/D BUFX2_99/A NOR2X1_15/A DFFSR_92/S
+ OAI22X1
XFILL_3_NOR2X1_32 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_13_DFFPOSX1_31 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_12_DFFSR_263 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_3_NAND3X1_35 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_4_OAI22X1_17 DFFSR_4/gnd DFFSR_98/S FILL
XDFFSR_153 INVX1_67/A CLKBUF1_2/Y BUFX2_67/Y DFFSR_201/S DFFSR_153/D INVX1_67/gnd
+ DFFSR_201/S DFFSR
XFILL_2_NAND2X1_108 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_51_6_0 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_3_OAI22X1_20 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_2_NAND3X1_38 BUFX2_98/A DFFSR_32/S FILL
XFILL_8_DFFSR_12 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_14_DFFSR_45 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_4_DFFSR_150 AND2X2_38/B DFFSR_23/S FILL
XFILL_1_BUFX2_80 BUFX2_79/A DFFSR_6/S FILL
XFILL_1_NAND3X1_41 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_2_OAI22X1_23 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_45_DFFSR_181 INVX1_3/gnd DFFSR_79/S FILL
XFILL_0_NAND3X1_44 BUFX2_99/A DFFSR_7/S FILL
XFILL_8_DFFSR_257 INVX1_39/gnd DFFSR_34/S FILL
XFILL_1_OAI22X1_26 INVX1_39/gnd DFFSR_54/S FILL
XFILL_35_DFFSR_184 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_23_DFFPOSX1_20 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_0_OAI22X1_29 INVX1_3/gnd DFFSR_79/S FILL
XFILL_25_DFFSR_187 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_49_DFFSR_62 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_15_DFFSR_190 INVX1_39/gnd DFFSR_34/S FILL
XFILL_7_NAND3X1_223 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_3_DFFPOSX1_42 INVX1_39/gnd DFFSR_34/S FILL
XINVX1_46 DFFSR_55/D DFFSR_4/gnd INVX1_46/Y DFFSR_4/S INVX1
XDFFSR_99 DFFSR_99/Q DFFSR_83/CLK DFFSR_73/R DFFSR_97/S DFFSR_91/Q XOR2X1_4/gnd DFFSR_97/S
+ DFFSR
XFILL_33_DFFSR_12 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_22_DFFSR_52 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_5_DFFSR_59 AND2X2_38/B DFFSR_59/S FILL
XFILL_11_DFFSR_92 BUFX2_99/A DFFSR_92/S FILL
XFILL_0_NOR2X1_69 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_48_DFFSR_108 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_38_DFFSR_111 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_8_NAND3X1_157 INVX1_3/gnd DFFSR_23/S FILL
XINVX1_164 INVX1_164/A BUFX2_8/gnd INVX1_164/Y DFFSR_81/S INVX1
XFILL_1_DFFSR_187 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_28_DFFSR_114 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_42_DFFSR_218 BUFX2_98/A DFFSR_32/S FILL
XFILL_1_NAND2X1_138 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_4_INVX1_161 INVX1_1/gnd DFFSR_53/S FILL
XFILL_7_AND2X2_28 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_18_DFFSR_117 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_32_DFFSR_221 AND2X2_38/B DFFSR_59/S FILL
XFILL_1_NAND2X1_8 INVX1_1/gnd DFFSR_53/S FILL
XFILL_22_DFFSR_224 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_41_DFFSR_19 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_2_INVX1_53 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_19_DFFSR_99 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_30_DFFSR_59 AND2X2_38/B DFFSR_59/S FILL
XFILL_12_DFFSR_227 BUFX2_7/gnd DFFSR_151/S FILL
XDFFSR_117 INVX1_37/A DFFSR_93/CLK DFFSR_5/R DFFSR_98/S DFFSR_109/Q BUFX2_77/gnd DFFSR_98/S
+ DFFSR
XFILL_22_DFFPOSX1_50 INVX1_1/gnd DFFSR_53/S FILL
XFILL_4_DFFSR_114 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_1_BUFX2_44 INVX1_3/gnd DFFSR_79/S FILL
XFILL_1_OAI22X1_7 AND2X2_38/B DFFSR_59/S FILL
XFILL_45_DFFSR_145 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_8_DFFSR_221 AND2X2_38/B DFFSR_59/S FILL
XFILL_35_DFFSR_148 INVX1_67/gnd DFFSR_175/S FILL
XFILL_8_DFFSR_2 BUFX2_79/A DFFSR_7/S FILL
XFILL_49_DFFSR_252 AND2X2_38/B DFFSR_23/S FILL
XFILL_25_DFFSR_151 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_39_DFFSR_255 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_38_DFFSR_66 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_49_DFFSR_26 BUFX2_79/A DFFSR_6/S FILL
XFILL_1_INVX1_198 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_7_NAND3X1_187 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_15_DFFSR_154 BUFX2_99/A DFFSR_7/S FILL
XFILL_29_DFFSR_258 DFFSR_5/gnd DFFSR_5/S FILL
XDFFSR_63 DFFSR_55/D CLKBUF1_38/Y DFFSR_15/R DFFSR_98/S DFFSR_63/D DFFSR_4/gnd DFFSR_98/S
+ DFFSR
XINVX1_10 DFFSR_50/Q BUFX2_77/gnd INVX1_10/Y DFFSR_5/S INVX1
XFILL_19_DFFSR_261 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_0_NAND2X1_168 BUFX2_79/A DFFSR_6/S FILL
XFILL_22_DFFSR_16 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_5_DFFSR_23 AND2X2_38/B DFFSR_23/S FILL
XFILL_11_DFFSR_56 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_0_NOR2X1_33 INVX1_3/gnd DFFSR_23/S FILL
XFILL_6_OR2X2_2 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_8_NAND3X1_121 INVX1_1/gnd DFFSR_97/S FILL
XINVX1_128 INVX1_62/A BUFX2_8/gnd INVX1_128/Y DFFSR_81/S INVX1
XFILL_4_NOR2X1_4 INVX1_1/gnd DFFSR_53/S FILL
XFILL_1_DFFSR_151 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_12_DFFPOSX1_25 BUFX2_79/A DFFSR_6/S FILL
XFILL_25_4_0 AND2X2_38/B DFFSR_23/S FILL
XFILL_32_DFFSR_6 BUFX2_79/A DFFSR_6/S FILL
XFILL_1_NAND2X1_102 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_42_DFFSR_182 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_4_INVX1_125 AND2X2_38/B DFFSR_59/S FILL
XFILL_46_DFFSR_73 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_5_DFFSR_258 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_32_DFFSR_185 INVX1_39/gnd DFFSR_54/S FILL
XFILL_23_6_1 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_22_DFFSR_188 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_2_DFFSR_70 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_2_INVX1_17 AND2X2_38/B DFFSR_59/S FILL
XFILL_5_5_0 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_19_DFFSR_63 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_30_DFFSR_23 AND2X2_38/B DFFSR_23/S FILL
XFILL_12_DFFSR_191 INVX1_67/gnd DFFSR_175/S FILL
XFILL_6_BUFX2_98 BUFX2_79/A DFFSR_7/S FILL
XFILL_22_DFFPOSX1_14 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_6_NAND3X1_217 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_45_DFFSR_109 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_2_DFFPOSX1_36 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_8_DFFSR_185 INVX1_39/gnd DFFSR_54/S FILL
XFILL_35_DFFSR_112 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_49_DFFSR_216 BUFX2_7/gnd DFFSR_216/S FILL
XAND2X2_32 BUFX2_58/Y AND2X2_34/B AND2X2_38/B AND2X2_32/Y DFFSR_23/S AND2X2
XFILL_25_DFFSR_115 INVX1_1/gnd DFFSR_97/S FILL
XFILL_39_DFFSR_219 INVX1_67/gnd DFFSR_175/S FILL
XFILL_27_DFFSR_70 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_38_DFFSR_30 BUFX2_98/A DFFSR_32/S FILL
XFILL_1_INVX1_162 INVX1_39/gnd DFFSR_34/S FILL
XFILL_4_AND2X2_29 AND2X2_38/B DFFSR_23/S FILL
XFILL_15_DFFSR_118 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_7_NAND3X1_151 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_29_DFFSR_222 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_19_DFFSR_225 INVX1_67/gnd DFFSR_175/S FILL
XFILL_0_NAND2X1_132 XOR2X1_1/gnd DFFSR_151/S FILL
XDFFSR_27 INVX1_22/A DFFSR_3/CLK DFFSR_3/R DFFSR_3/S DFFSR_3/Q DFFSR_28/gnd DFFSR_3/S
+ DFFSR
XFILL_11_DFFSR_20 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_8_OAI22X1_5 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_2_NOR3X1_1 INVX1_3/gnd DFFSR_79/S FILL
XFILL_17_4 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_1_DFFSR_115 INVX1_1/gnd DFFSR_97/S FILL
XFILL_21_DFFPOSX1_44 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_42_DFFSR_146 BUFX2_79/A DFFSR_7/S FILL
XFILL_33_1_1 INVX1_1/gnd DFFSR_53/S FILL
XFILL_46_DFFSR_37 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_35_DFFSR_77 BUFX2_98/A DFFSR_32/S FILL
XFILL_5_DFFSR_222 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_32_DFFSR_149 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_46_DFFSR_253 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_5_NAND3X1_247 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_22_DFFSR_152 INVX1_1/gnd DFFSR_53/S FILL
XFILL_31_3_2 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_2_DFFSR_34 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_19_DFFSR_27 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_36_DFFSR_256 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_12_DFFSR_155 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_6_BUFX2_62 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_26_DFFSR_259 BUFX2_79/A DFFSR_6/S FILL
XFILL_8_OAI21X1_103 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_16_DFFSR_262 BUFX2_98/A DFFSR_32/S FILL
XFILL_20_CLKBUF1_17 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_6_NAND3X1_181 INVX1_39/gnd DFFSR_54/S FILL
XFILL_43_DFFSR_84 BUFX2_99/A DFFSR_7/S FILL
XFILL_19_CLKBUF1_20 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_8_DFFSR_149 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_18_CLKBUF1_23 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_49_DFFSR_180 DFFSR_34/gnd DFFSR_34/S FILL
XNAND3X1_217 AOI21X1_25/Y NAND3X1_217/B NAND3X1_216/Y DFFSR_46/gnd NAND2X1_99/A DFFSR_54/S
+ NAND3X1
XFILL_39_DFFSR_183 INVX1_67/gnd DFFSR_175/S FILL
XFILL_17_CLKBUF1_26 INVX1_1/gnd DFFSR_53/S FILL
XFILL_1_INVX1_126 INVX1_3/gnd DFFSR_23/S FILL
XFILL_27_DFFSR_34 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_16_DFFSR_74 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_2_DFFSR_259 BUFX2_79/A DFFSR_6/S FILL
XFILL_7_NAND3X1_115 BUFX2_79/A DFFSR_7/S FILL
XFILL_3_BUFX2_1 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_29_DFFSR_186 BUFX2_99/A DFFSR_92/S FILL
XFILL_16_CLKBUF1_29 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_11_DFFPOSX1_19 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_19_DFFSR_189 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_15_CLKBUF1_32 DFFSR_1/gnd DFFSR_81/S FILL
XNOR2X1_71 NOR2X1_70/B NOR2X1_71/B INVX1_1/gnd NOR2X1_71/Y DFFSR_97/S NOR2X1
XFILL_14_CLKBUF1_35 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_13_CLKBUF1_38 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_4_NOR2X1_68 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_12_CLKBUF1_41 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_42_DFFSR_110 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_7_DFFSR_88 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_35_DFFSR_41 BUFX2_98/A DFFSR_6/S FILL
XFILL_11_CLKBUF1_44 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_24_DFFSR_81 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_5_DFFSR_186 BUFX2_99/A DFFSR_92/S FILL
XFILL_32_DFFSR_113 BUFX2_99/A DFFSR_92/S FILL
XFILL_46_DFFSR_217 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_10_CLKBUF1_47 BUFX2_98/A DFFSR_32/S FILL
XFILL_5_NAND3X1_211 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_22_DFFSR_116 INVX1_3/gnd DFFSR_23/S FILL
XFILL_36_DFFSR_220 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_1_DFFPOSX1_30 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_1_AND2X2_30 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_12_DFFSR_119 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_6_BUFX2_26 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_5_NAND2X1_7 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_26_DFFSR_223 INVX1_39/gnd DFFSR_34/S FILL
XFILL_16_DFFSR_226 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_16_NOR3X1_5 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_44_DFFSR_9 BUFX2_79/A DFFSR_6/S FILL
XFILL_6_NAND3X1_145 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_10_DFFPOSX1_49 BUFX2_99/A DFFSR_92/S FILL
XFILL_4_INVX1_82 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_43_DFFSR_48 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_32_DFFSR_88 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_8_DFFSR_113 BUFX2_99/A DFFSR_92/S FILL
XFILL_5_OAI22X1_6 BUFX2_98/A DFFSR_32/S FILL
XFILL_49_DFFSR_144 DFFSR_46/gnd DFFSR_62/S FILL
XNAND3X1_181 INVX1_158/A OAI21X1_47/Y NAND2X1_83/Y INVX1_39/gnd AOI22X1_24/A DFFSR_54/S
+ NAND3X1
XFILL_39_DFFSR_147 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_16_DFFSR_38 BUFX2_98/A DFFSR_6/S FILL
XFILL_2_DFFSR_223 INVX1_39/gnd DFFSR_34/S FILL
XFILL_39_4 BUFX2_79/A DFFSR_7/S FILL
XFILL_3_BUFX2_73 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_29_DFFSR_150 AND2X2_38/B DFFSR_23/S FILL
XFILL_43_DFFSR_254 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_20_DFFPOSX1_38 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_19_DFFSR_153 INVX1_67/gnd DFFSR_201/S FILL
XFILL_33_DFFSR_257 INVX1_39/gnd DFFSR_34/S FILL
XNOR2X1_35 NOR2X1_35/A OAI21X1_9/Y OR2X2_2/gnd NOR2X1_35/Y DFFSR_216/S NOR2X1
XFILL_4_NAND3X1_241 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_23_DFFSR_260 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_40_DFFSR_95 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_4_NOR2X1_32 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_13_DFFSR_263 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_1_AND2X2_4 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_7_DFFSR_52 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_13_DFFSR_85 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_24_DFFSR_45 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_5_DFFSR_150 AND2X2_38/B DFFSR_23/S FILL
XFILL_46_DFFSR_181 INVX1_3/gnd DFFSR_79/S FILL
XFILL_10_CLKBUF1_11 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_5_NAND3X1_175 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_9_DFFSR_257 INVX1_39/gnd DFFSR_34/S FILL
XFILL_36_DFFSR_184 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_26_DFFSR_187 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_9_CLKBUF1_14 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_10_DFFSR_7 BUFX2_79/A DFFSR_7/S FILL
XFILL_8_CLKBUF1_17 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_16_DFFSR_190 INVX1_39/gnd DFFSR_34/S FILL
XFILL_6_NAND3X1_109 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_32_4_0 INVX1_1/gnd DFFSR_97/S FILL
XFILL_7_CLKBUF1_20 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_10_DFFPOSX1_13 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_43_DFFSR_12 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_32_DFFSR_52 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_4_INVX1_46 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_4_DFFSR_99 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_21_DFFSR_92 BUFX2_99/A DFFSR_92/S FILL
XFILL_6_CLKBUF1_23 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_1_NOR2X1_69 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_49_DFFSR_108 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_5_CLKBUF1_26 INVX1_1/gnd DFFSR_53/S FILL
XFILL_30_6_1 XOR2X1_4/gnd DFFSR_91/S FILL
XNAND3X1_145 AOI21X1_12/B AOI21X1_12/C AOI21X1_12/A DFFSR_1/gnd AOI22X1_20/A DFFSR_81/S
+ NAND3X1
XFILL_39_DFFSR_111 DFFSR_8/gnd DFFSR_8/S FILL
XCLKBUF1_23 BUFX2_2/Y DFFSR_4/gnd DFFSR_85/CLK DFFSR_98/S CLKBUF1
XOR2X2_3 OR2X2_3/A OR2X2_3/B OR2X2_3/gnd OR2X2_3/Y DFFSR_4/S OR2X2
XFILL_4_CLKBUF1_29 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_2_DFFSR_187 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_3_BUFX2_37 INVX1_1/gnd DFFSR_97/S FILL
XFILL_29_DFFSR_114 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_43_DFFSR_218 BUFX2_98/A DFFSR_32/S FILL
XFILL_3_CLKBUF1_32 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_8_AND2X2_28 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_19_DFFSR_117 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_2_CLKBUF1_35 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_33_DFFSR_221 AND2X2_38/B DFFSR_59/S FILL
XFILL_31_DFFSR_3 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_2_NAND2X1_8 INVX1_1/gnd DFFSR_53/S FILL
XFILL_23_DFFSR_224 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_1_CLKBUF1_38 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_4_NAND3X1_205 INVX1_1/gnd DFFSR_53/S FILL
XFILL_29_DFFSR_99 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_1_INVX1_93 INVX1_3/gnd DFFSR_23/S FILL
XFILL_40_DFFSR_59 AND2X2_38/B DFFSR_59/S FILL
XFILL_13_DFFSR_227 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_0_DFFPOSX1_24 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_0_CLKBUF1_41 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_7_DFFSR_16 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_13_DFFSR_49 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_5_DFFSR_114 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_0_BUFX2_84 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_2_OAI22X1_7 AND2X2_38/B DFFSR_59/S FILL
XFILL_46_DFFSR_145 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_5_NAND3X1_139 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_9_DFFSR_221 AND2X2_38/B DFFSR_59/S FILL
XFILL_36_DFFSR_148 INVX1_67/gnd DFFSR_175/S FILL
XFILL_50_DFFSR_252 AND2X2_38/B DFFSR_23/S FILL
XFILL_26_DFFSR_151 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_48_DFFSR_66 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_40_DFFSR_255 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_2_INVX1_198 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_16_DFFSR_154 BUFX2_99/A DFFSR_7/S FILL
XFILL_30_DFFSR_258 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_20_DFFSR_261 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_32_DFFSR_16 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_4_DFFSR_63 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_19_DFFPOSX1_32 INVX1_67/gnd DFFSR_201/S FILL
XFILL_21_DFFSR_56 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_10_DFFSR_96 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_40_1_1 BUFX2_98/A DFFSR_6/S FILL
XFILL_1_NOR2X1_33 INVX1_3/gnd DFFSR_23/S FILL
XFILL_10_DFFSR_264 DFFSR_4/gnd DFFSR_98/S FILL
XNAND3X1_109 DFFSR_198/D BUFX2_34/Y BUFX2_23/Y XOR2X1_1/gnd NAND3X1_111/A DFFSR_151/S
+ NAND3X1
XFILL_3_NAND3X1_235 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_38_3_2 BUFX2_79/A DFFSR_7/S FILL
XFILL_2_DFFSR_151 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_43_DFFSR_182 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_6_DFFSR_258 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_33_DFFSR_185 INVX1_39/gnd DFFSR_54/S FILL
XFILL_23_DFFSR_188 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_4_NAND3X1_169 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_29_DFFSR_63 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_1_INVX1_57 BUFX2_98/A DFFSR_32/S FILL
XFILL_40_DFFSR_23 AND2X2_38/B DFFSR_23/S FILL
XFILL_13_DFFSR_191 INVX1_67/gnd DFFSR_175/S FILL
XFILL_9_DFFPOSX1_43 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_13_DFFSR_13 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_0_BUFX2_48 AND2X2_38/B DFFSR_59/S FILL
XFILL_46_DFFSR_109 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_5_NAND3X1_103 AND2X2_38/B DFFSR_23/S FILL
XFILL_9_DFFSR_185 INVX1_39/gnd DFFSR_54/S FILL
XFILL_36_DFFSR_112 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_50_DFFSR_216 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_26_DFFSR_115 INVX1_1/gnd DFFSR_97/S FILL
XFILL_40_DFFSR_219 INVX1_67/gnd DFFSR_175/S FILL
XFILL_48_DFFSR_30 BUFX2_98/A DFFSR_32/S FILL
XFILL_2_INVX1_162 INVX1_39/gnd DFFSR_34/S FILL
XFILL_37_DFFSR_70 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_5_AND2X2_29 AND2X2_38/B DFFSR_23/S FILL
XFILL_16_DFFSR_118 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_30_DFFSR_222 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_20_DFFSR_225 INVX1_67/gnd DFFSR_175/S FILL
XFILL_4_DFFSR_27 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_10_DFFSR_60 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_21_DFFSR_20 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_10_DFFSR_228 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_3_NAND3X1_199 INVX1_1/gnd DFFSR_97/S FILL
XFILL_9_OAI22X1_5 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_3_NOR2X1_8 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_2_DFFSR_115 INVX1_1/gnd DFFSR_97/S FILL
XFILL_43_DFFSR_146 BUFX2_79/A DFFSR_7/S FILL
XFILL_45_DFFSR_77 BUFX2_98/A DFFSR_32/S FILL
XFILL_6_DFFSR_222 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_33_DFFSR_149 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_47_DFFSR_253 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_23_DFFSR_152 INVX1_1/gnd DFFSR_53/S FILL
XFILL_4_NAND3X1_133 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_29_DFFSR_27 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_37_DFFSR_256 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_1_DFFSR_74 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_1_INVX1_21 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_18_DFFSR_67 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_13_DFFSR_155 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_27_DFFSR_259 BUFX2_79/A DFFSR_6/S FILL
XFILL_6_NAND2X1_169 INVX1_1/gnd DFFSR_53/S FILL
XFILL_17_DFFSR_262 BUFX2_98/A DFFSR_32/S FILL
XFILL_0_BUFX2_12 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_5_XOR2X1_4 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_21_DFFPOSX1_2 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_9_DFFSR_149 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_43_DFFSR_6 BUFX2_79/A DFFSR_6/S FILL
XFILL_20_DFFPOSX1_5 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_18_DFFPOSX1_26 AND2X2_38/B DFFSR_23/S FILL
XFILL_50_DFFSR_180 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_19_DFFPOSX1_8 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_12_1_2 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_40_DFFSR_183 INVX1_67/gnd DFFSR_175/S FILL
XFILL_2_INVX1_126 INVX1_3/gnd DFFSR_23/S FILL
XFILL_9_DFFSR_81 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_26_DFFSR_74 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_37_DFFSR_34 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_2_NAND3X1_229 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_3_DFFSR_259 BUFX2_79/A DFFSR_6/S FILL
XFILL_30_DFFSR_186 BUFX2_99/A DFFSR_92/S FILL
XFILL_20_DFFSR_189 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_10_DFFSR_24 BUFX2_98/A DFFSR_6/S FILL
XFILL_10_DFFSR_192 INVX1_1/gnd DFFSR_97/S FILL
XFILL_5_NOR2X1_68 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_3_NAND3X1_163 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_1_NOR3X1_5 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_8_DFFPOSX1_37 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_43_DFFSR_110 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_45_DFFSR_41 BUFX2_98/A DFFSR_6/S FILL
XFILL_34_DFFSR_81 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_6_DFFSR_186 BUFX2_99/A DFFSR_92/S FILL
XFILL_33_DFFSR_113 BUFX2_99/A DFFSR_92/S FILL
XFILL_47_DFFSR_217 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_23_DFFSR_116 INVX1_3/gnd DFFSR_23/S FILL
XFILL_37_DFFSR_220 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_1_DFFSR_38 BUFX2_98/A DFFSR_6/S FILL
XFILL_18_DFFSR_31 BUFX2_79/A DFFSR_6/S FILL
XFILL_39_4_0 BUFX2_79/A DFFSR_6/S FILL
XFILL_2_AND2X2_30 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_13_DFFSR_119 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_6_NAND2X1_7 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_5_BUFX2_66 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_27_DFFSR_223 INVX1_39/gnd DFFSR_34/S FILL
XFILL_6_NAND2X1_133 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_17_DFFSR_226 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_37_6_1 BUFX2_99/A DFFSR_7/S FILL
XXOR2X1_8 XOR2X1_8/A XOR2X1_8/B OR2X2_4/gnd OR2X2_4/B DFFSR_3/S XOR2X1
XFILL_11_XOR2X1_1 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_42_DFFSR_88 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_9_DFFSR_113 BUFX2_99/A DFFSR_92/S FILL
XNAND2X1_169 DFFSR_91/S DFFPOSX1_5/Q INVX1_1/gnd AOI21X1_60/B DFFSR_53/S NAND2X1
XFILL_6_OAI22X1_6 BUFX2_98/A DFFSR_32/S FILL
XFILL_50_DFFSR_144 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_4_OAI21X1_115 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_8_AOI21X1_61 AND2X2_38/B DFFSR_59/S FILL
XFILL_27_DFFPOSX1_45 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_40_DFFSR_147 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_9_DFFSR_45 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_15_DFFSR_78 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_26_DFFSR_38 BUFX2_98/A DFFSR_6/S FILL
XFILL_7_AOI21X1_64 AND2X2_38/B DFFSR_59/S FILL
XFILL_3_DFFSR_223 INVX1_39/gnd DFFSR_34/S FILL
XFILL_2_NAND3X1_193 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_43_1 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_30_DFFSR_150 AND2X2_38/B DFFSR_23/S FILL
XFILL_6_AOI21X1_67 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_44_DFFSR_254 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_20_DFFSR_153 INVX1_67/gnd DFFSR_201/S FILL
XFILL_5_AOI21X1_70 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_34_DFFSR_257 INVX1_39/gnd DFFSR_34/S FILL
XFILL_10_DFFSR_156 OR2X2_2/gnd DFFSR_175/S FILL
XAOI21X1_67 AOI21X1_67/A XOR2X1_13/Y AOI21X1_67/C NOR3X1_6/gnd AOI21X1_67/Y DFFSR_91/S
+ AOI21X1
XFILL_24_DFFSR_260 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_50_DFFSR_95 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_5_NOR2X1_32 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_3_NAND3X1_127 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_14_DFFSR_263 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_5_NAND2X1_163 INVX1_67/gnd DFFSR_201/S FILL
XFILL_34_DFFSR_45 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_6_DFFSR_92 BUFX2_99/A DFFSR_92/S FILL
XFILL_23_DFFSR_85 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_6_DFFSR_150 AND2X2_38/B DFFSR_23/S FILL
XFILL_47_DFFSR_181 INVX1_3/gnd DFFSR_79/S FILL
XFILL_37_DFFSR_184 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_0_DFFSR_260 BUFX2_77/gnd DFFSR_5/S FILL
XBUFX2_70 BUFX2_60/A BUFX2_77/gnd BUFX2_70/Y DFFSR_5/S BUFX2
XFILL_47_1_1 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_5_BUFX2_30 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_17_DFFPOSX1_20 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_27_DFFSR_187 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_17_DFFSR_190 INVX1_39/gnd DFFSR_34/S FILL
XFILL_1_NAND3X1_223 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_9_DFFPOSX1_2 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_45_3_2 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_8_DFFPOSX1_5 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_42_DFFSR_52 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_31_DFFSR_92 BUFX2_99/A DFFSR_92/S FILL
XFILL_3_INVX1_86 DFFSR_46/gnd DFFSR_54/S FILL
XNAND2X1_133 DFFSR_175/S DFFSR_266/Q BUFX2_72/gnd NAND2X1_133/Y DFFSR_201/S NAND2X1
XFILL_2_NOR2X1_69 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_50_DFFSR_108 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_7_DFFPOSX1_8 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_8_AOI21X1_25 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_40_DFFSR_111 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_15_DFFSR_42 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_7_AOI21X1_28 AND2X2_38/B DFFSR_23/S FILL
XFILL_2_NAND3X1_157 INVX1_3/gnd DFFSR_23/S FILL
XFILL_3_DFFSR_187 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_2_BUFX2_77 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_30_DFFSR_114 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_6_AOI21X1_31 INVX1_39/gnd DFFSR_34/S FILL
XFILL_44_DFFSR_218 BUFX2_98/A DFFSR_32/S FILL
XFILL_9_AND2X2_28 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_20_DFFSR_117 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_7_DFFPOSX1_31 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_5_AOI21X1_34 INVX1_39/gnd DFFSR_34/S FILL
XFILL_34_DFFSR_221 AND2X2_38/B DFFSR_59/S FILL
XFILL_10_DFFSR_120 INVX1_3/gnd DFFSR_23/S FILL
XAOI21X1_31 AOI21X1_22/C AOI21X1_22/B OAI21X1_73/A INVX1_39/gnd AOI21X1_31/Y DFFSR_34/S
+ AOI21X1
XFILL_4_AOI21X1_37 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_3_NAND2X1_8 INVX1_1/gnd DFFSR_53/S FILL
XFILL_13_2_0 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_24_DFFSR_224 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_39_DFFSR_99 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_50_DFFSR_59 AND2X2_38/B DFFSR_59/S FILL
XFILL_14_DFFSR_227 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_3_AOI21X1_40 INVX1_39/gnd DFFSR_54/S FILL
XFILL_16_DFFPOSX1_50 INVX1_1/gnd DFFSR_53/S FILL
XFILL_2_AOI21X1_43 INVX1_3/gnd DFFSR_79/S FILL
XFILL_11_4_1 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_0_AND2X2_8 BUFX2_99/A DFFSR_7/S FILL
XFILL_6_DFFSR_56 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_23_DFFSR_49 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_5_NAND2X1_127 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_1_AOI21X1_46 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_6_DFFSR_114 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_12_DFFSR_89 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_3_OAI22X1_7 AND2X2_38/B DFFSR_59/S FILL
XFILL_47_DFFSR_145 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_0_AOI21X1_49 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_37_DFFSR_148 INVX1_67/gnd DFFSR_175/S FILL
XFILL_0_DFFSR_224 BUFX2_7/gnd DFFSR_151/S FILL
XBUFX2_34 BUFX2_34/A DFFSR_46/gnd BUFX2_34/Y DFFSR_54/S BUFX2
XFILL_27_DFFSR_151 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_3_OAI21X1_109 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_26_DFFPOSX1_39 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_41_DFFSR_255 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_3_INVX1_198 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_48_6 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_17_DFFSR_154 BUFX2_99/A DFFSR_7/S FILL
XFILL_8_OAI21X1_73 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_1_NAND3X1_187 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_31_DFFSR_258 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_21_DFFSR_261 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_6_NAND2X1_94 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_7_OAI21X1_76 INVX1_1/gnd DFFSR_53/S FILL
XFILL_42_DFFSR_16 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_31_DFFSR_56 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_20_DFFSR_96 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_3_INVX1_50 BUFX2_98/A DFFSR_6/S FILL
XFILL_2_NOR2X1_33 INVX1_3/gnd DFFSR_23/S FILL
XFILL_6_OAI21X1_79 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_5_NAND2X1_97 INVX1_1/gnd DFFSR_97/S FILL
XFILL_11_DFFSR_264 DFFSR_4/gnd DFFSR_98/S FILL
XNAND2X1_94 NOR2X1_69/Y XOR2X1_4/Y OR2X2_6/gnd AOI22X1_26/A DFFSR_92/S NAND2X1
XFILL_5_OAI21X1_82 DFFSR_28/gnd DFFSR_8/S FILL
XOAI21X1_79 INVX1_175/Y INVX1_161/Y INVX1_176/Y DFFSR_8/gnd OAI21X1_79/Y DFFSR_8/S
+ OAI21X1
XFILL_3_DFFSR_151 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_2_NAND3X1_121 INVX1_1/gnd DFFSR_97/S FILL
XFILL_2_BUFX2_41 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_4_OAI21X1_85 INVX1_39/gnd DFFSR_54/S FILL
XFILL_44_DFFSR_182 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_3_OAI21X1_88 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_7_DFFSR_258 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_4_NAND2X1_157 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_34_DFFSR_185 INVX1_39/gnd DFFSR_54/S FILL
XFILL_2_OAI21X1_91 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_21_DFFSR_7 BUFX2_79/A DFFSR_7/S FILL
XFILL_24_DFFSR_188 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_1_OAI21X1_94 INVX1_67/gnd DFFSR_175/S FILL
XFILL_39_DFFSR_63 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_50_DFFSR_23 AND2X2_38/B DFFSR_23/S FILL
XFILL_0_INVX1_97 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_14_DFFSR_191 INVX1_67/gnd DFFSR_175/S FILL
XFILL_0_OAI21X1_97 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_16_DFFPOSX1_14 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_6_DFFSR_20 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_23_DFFSR_13 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_19_1_2 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_12_DFFSR_53 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_5_BUFX2_8 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_1_AOI21X1_10 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_47_DFFSR_109 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_0_NAND3X1_217 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_0_AOI21X1_13 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_1_0_1 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_37_DFFSR_112 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_5_NOR2X1_1 BUFX2_99/A DFFSR_92/S FILL
XFILL_0_DFFSR_188 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_27_DFFSR_115 INVX1_1/gnd DFFSR_97/S FILL
XFILL_42_DFFSR_3 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_41_DFFSR_219 INVX1_67/gnd DFFSR_175/S FILL
XFILL_3_INVX1_162 INVX1_39/gnd DFFSR_34/S FILL
XFILL_47_DFFSR_70 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_6_AND2X2_29 AND2X2_38/B DFFSR_23/S FILL
XFILL_17_DFFSR_118 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_8_OAI21X1_37 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_31_DFFSR_222 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_1_NAND3X1_151 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_0_NAND2X1_9 BUFX2_79/A DFFSR_6/S FILL
XFILL_21_DFFSR_225 INVX1_67/gnd DFFSR_175/S FILL
XFILL_6_NAND2X1_58 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_7_OAI21X1_40 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_3_INVX1_14 BUFX2_98/A DFFSR_6/S FILL
XFILL_20_DFFSR_60 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_31_DFFSR_20 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_3_DFFSR_67 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_6_DFFPOSX1_25 BUFX2_79/A DFFSR_6/S FILL
XFILL_5_NAND2X1_61 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_6_OAI21X1_43 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_11_DFFSR_228 XOR2X1_1/gnd DFFSR_208/S FILL
XNAND2X1_58 BUFX2_56/Y INVX1_133/A BUFX2_8/gnd XOR2X1_1/B DFFSR_81/S NAND2X1
XFILL_5_OAI21X1_46 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_4_NAND2X1_64 DFFSR_46/gnd DFFSR_62/S FILL
XOAI21X1_43 AOI21X1_16/Y AOI21X1_17/Y INVX1_155/A BUFX2_7/gnd OAI21X1_43/Y DFFSR_151/S
+ OAI21X1
XFILL_3_DFFSR_115 INVX1_1/gnd DFFSR_97/S FILL
XFILL_3_NAND2X1_67 AND2X2_38/B DFFSR_59/S FILL
XFILL_46_4_0 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_4_OAI21X1_49 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_0_OAI22X1_8 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_44_DFFSR_146 BUFX2_79/A DFFSR_7/S FILL
XFILL_15_DFFPOSX1_44 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_2_NAND2X1_70 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_3_OAI21X1_52 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_7_DFFSR_222 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_4_NAND2X1_121 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_34_DFFSR_149 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_1_NAND2X1_73 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_2_OAI21X1_55 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_44_6_1 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_48_DFFSR_253 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_24_DFFSR_152 INVX1_1/gnd DFFSR_53/S FILL
XFILL_0_NAND2X1_76 INVX1_3/gnd DFFSR_23/S FILL
XFILL_1_OAI21X1_58 INVX1_39/gnd DFFSR_54/S FILL
XFILL_39_DFFSR_27 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_38_DFFSR_256 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_0_INVX1_61 INVX1_39/gnd DFFSR_54/S FILL
XFILL_10_AOI22X1_24 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_0_INVX1_199 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_28_DFFSR_67 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_14_DFFSR_155 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_28_DFFSR_259 BUFX2_79/A DFFSR_6/S FILL
XFILL_0_OAI21X1_61 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_2_OAI21X1_103 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_18_DFFSR_262 BUFX2_98/A DFFSR_32/S FILL
XFILL_25_DFFPOSX1_33 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_9_AOI22X1_27 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_12_DFFSR_17 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_0_NAND3X1_181 INVX1_39/gnd DFFSR_54/S FILL
XNOR2X1_5 NOR3X1_2/C NOR2X1_5/B OR2X2_6/gnd NOR2X1_5/Y DFFSR_53/S NOR2X1
XFILL_0_DFFSR_152 INVX1_1/gnd DFFSR_53/S FILL
XDFFSR_262 DFFSR_6/D DFFSR_2/CLK DFFSR_257/R DFFSR_32/S DFFSR_262/D BUFX2_98/A DFFSR_32/S
+ DFFSR
XFILL_41_DFFSR_183 INVX1_67/gnd DFFSR_175/S FILL
XFILL_3_INVX1_126 INVX1_3/gnd DFFSR_23/S FILL
XFILL_36_DFFSR_74 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_47_DFFSR_34 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_4_DFFSR_259 BUFX2_79/A DFFSR_6/S FILL
XFILL_1_NAND3X1_115 BUFX2_79/A DFFSR_7/S FILL
XFILL_31_DFFSR_186 BUFX2_99/A DFFSR_92/S FILL
XFILL_6_NAND2X1_22 BUFX2_99/A DFFSR_7/S FILL
XFILL_21_DFFSR_189 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_20_DFFSR_24 BUFX2_98/A DFFSR_6/S FILL
XFILL_3_DFFSR_31 BUFX2_79/A DFFSR_6/S FILL
XFILL_5_NAND2X1_25 BUFX2_99/A DFFSR_7/S FILL
XFILL_11_DFFSR_192 INVX1_1/gnd DFFSR_97/S FILL
XFILL_3_NAND2X1_151 DFFSR_1/gnd DFFSR_81/S FILL
XNAND2X1_22 DFFSR_46/D AND2X2_5/Y BUFX2_99/A NAND2X1_22/Y DFFSR_7/S NAND2X1
XFILL_5_OAI21X1_10 BUFX2_79/A DFFSR_7/S FILL
XFILL_4_NAND2X1_28 AND2X2_38/B DFFSR_59/S FILL
XFILL_6_NOR2X1_68 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_8_2 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_3_NAND2X1_31 INVX1_3/gnd DFFSR_23/S FILL
XFILL_4_OAI21X1_13 INVX1_39/gnd DFFSR_54/S FILL
XFILL_9_DFFSR_6 BUFX2_79/A DFFSR_6/S FILL
XDFFPOSX1_25 NAND2X1_167/B CLKBUF1_46/Y AOI21X1_60/Y BUFX2_79/A DFFSR_6/S DFFPOSX1
XFILL_44_DFFSR_110 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_54_1_1 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_3_OAI21X1_16 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_2_NAND2X1_34 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_44_DFFSR_81 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_7_DFFSR_186 BUFX2_99/A DFFSR_92/S FILL
XFILL_34_DFFSR_113 BUFX2_99/A DFFSR_92/S FILL
XFILL_1_NAND2X1_37 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_2_OAI21X1_19 BUFX2_98/A DFFSR_32/S FILL
XFILL_48_DFFSR_217 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_24_DFFSR_116 INVX1_3/gnd DFFSR_23/S FILL
XFILL_8_NAND3X1_93 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_52_3_2 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_0_NAND2X1_40 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_1_OAI21X1_22 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_38_DFFSR_220 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_0_INVX1_25 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_0_DFFSR_78 OR2X2_3/gnd DFFSR_4/S FILL
XAOI21X1_1 AOI21X1_1/A AOI21X1_1/B AOI21X1_1/C DFFSR_34/gnd AOI21X1_1/Y DFFSR_34/S
+ AOI21X1
XFILL_0_INVX1_163 INVX1_39/gnd DFFSR_54/S FILL
XFILL_3_AND2X2_30 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_28_DFFSR_31 BUFX2_79/A DFFSR_6/S FILL
XFILL_17_DFFSR_71 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_14_DFFSR_119 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_7_NAND3X1_96 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_28_DFFSR_223 INVX1_39/gnd DFFSR_34/S FILL
XFILL_0_OAI21X1_25 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_6_NAND3X1_99 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_18_DFFSR_226 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_7_OR2X2_6 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_4_XOR2X1_8 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_0_NAND3X1_145 DFFSR_1/gnd DFFSR_81/S FILL
XNAND3X1_99 BUFX2_94/A AND2X2_16/Y BUFX2_32/Y OR2X2_1/gnd AND2X2_23/A DFFSR_51/S NAND3X1
XFILL_7_OAI22X1_6 BUFX2_98/A DFFSR_32/S FILL
XFILL_5_DFFPOSX1_19 DFFSR_34/gnd DFFSR_1/S FILL
XDFFSR_226 DFFSR_234/D DFFSR_5/CLK BUFX2_65/Y DFFSR_98/S DFFSR_218/Q DFFSR_4/gnd DFFSR_98/S
+ DFFSR
XFILL_0_DFFSR_116 INVX1_3/gnd DFFSR_23/S FILL
XFILL_2_NAND2X1_181 BUFX2_99/A DFFSR_92/S FILL
XFILL_30_3 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_20_2_0 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_41_DFFSR_147 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_8_DFFSR_85 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_25_DFFSR_78 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_36_DFFSR_38 BUFX2_98/A DFFSR_6/S FILL
XFILL_4_DFFSR_223 INVX1_39/gnd DFFSR_34/S FILL
XFILL_31_DFFSR_150 AND2X2_38/B DFFSR_23/S FILL
XFILL_45_DFFSR_254 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_21_DFFSR_153 INVX1_67/gnd DFFSR_201/S FILL
XFILL_14_DFFPOSX1_38 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_18_4_1 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_35_DFFSR_257 INVX1_39/gnd DFFSR_34/S FILL
XFILL_11_DFFSR_156 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_3_NAND2X1_115 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_25_DFFSR_260 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_0_3_0 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_2_AOI22X1_12 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_6_NOR2X1_32 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_15_DFFSR_263 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_11_OAI22X1_33 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_16_6_2 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_1_AOI22X1_15 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_17_NOR3X1_2 INVX1_1/gnd DFFSR_53/S FILL
XFILL_10_OAI22X1_36 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_0_AOI22X1_18 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_44_DFFSR_45 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_33_DFFSR_85 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_7_DFFSR_150 AND2X2_38/B DFFSR_23/S FILL
XFILL_24_DFFPOSX1_27 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_48_DFFSR_181 INVX1_3/gnd DFFSR_79/S FILL
XFILL_8_NAND3X1_57 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_9_OAI22X1_39 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_8_NAND3X1_230 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_0_DFFSR_42 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_38_DFFSR_184 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_0_INVX1_127 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_17_DFFSR_35 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_7_NAND3X1_60 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_1_DFFSR_260 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_4_BUFX2_70 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_8_OAI22X1_42 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_4_DFFPOSX1_49 BUFX2_99/A DFFSR_92/S FILL
XFILL_28_DFFSR_187 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_7_OAI22X1_45 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_6_NAND3X1_63 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_18_DFFSR_190 INVX1_39/gnd DFFSR_34/S FILL
XFILL_5_NAND3X1_66 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_6_OAI22X1_48 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_0_NAND3X1_109 XOR2X1_1/gnd DFFSR_151/S FILL
XNAND3X1_63 NAND3X1_61/Y NAND3X1_63/B AOI22X1_8/Y DFFSR_28/gnd NOR2X1_29/B DFFSR_3/S
+ NAND3X1
XFILL_10_XOR2X1_5 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_4_NAND3X1_69 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_9_NAND3X1_164 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_5_OAI22X1_51 INVX1_39/gnd DFFSR_54/S FILL
XFILL_41_DFFSR_92 BUFX2_99/A DFFSR_92/S FILL
XFILL_3_NOR2X1_69 OR2X2_6/gnd DFFSR_92/S FILL
XOAI22X1_48 INVX1_115/Y OAI22X1_45/B INVX1_116/Y OAI22X1_45/D XOR2X1_4/gnd NOR2X1_57/A
+ DFFSR_91/S OAI22X1
XFILL_51_DFFSR_108 OR2X2_6/gnd DFFSR_92/S FILL
XDFFSR_190 INVX1_98/A CLKBUF1_17/Y BUFX2_69/Y DFFSR_34/S DFFSR_190/D INVX1_39/gnd
+ DFFSR_34/S DFFSR
XFILL_3_NAND3X1_72 INVX1_39/gnd DFFSR_34/S FILL
XFILL_2_NAND2X1_145 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_2_AND2X2_1 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_41_DFFSR_111 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_2_NAND3X1_75 BUFX2_79/A DFFSR_7/S FILL
XFILL_25_DFFSR_42 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_8_DFFSR_49 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_14_DFFSR_82 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_4_DFFSR_187 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_31_DFFSR_114 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_1_NAND3X1_78 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_45_DFFSR_218 BUFX2_98/A DFFSR_32/S FILL
XFILL_21_DFFSR_117 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_0_NAND3X1_81 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_35_DFFSR_221 AND2X2_38/B DFFSR_59/S FILL
XFILL_0_AND2X2_31 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_26_1_2 INVX1_3/gnd DFFSR_23/S FILL
XFILL_11_DFFSR_120 INVX1_3/gnd DFFSR_23/S FILL
XFILL_4_NAND2X1_8 INVX1_1/gnd DFFSR_53/S FILL
XFILL_25_DFFSR_224 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_49_DFFSR_99 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_20_DFFSR_4 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_8_0_1 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_15_DFFSR_227 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_5_DFFSR_96 DFFSR_4/gnd DFFSR_4/S FILL
XINVX1_83 INVX1_83/A INVX1_39/gnd INVX1_83/Y DFFSR_54/S INVX1
XFILL_33_DFFSR_49 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_7_DFFSR_114 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_22_DFFSR_89 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_6_2_2 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_9_NAND3X1_18 BUFX2_79/A DFFSR_7/S FILL
XFILL_4_OAI22X1_7 AND2X2_38/B DFFSR_59/S FILL
XFILL_48_DFFSR_145 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_8_NAND3X1_21 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_4_BUFX2_5 AND2X2_38/B DFFSR_59/S FILL
XFILL_38_DFFSR_148 INVX1_67/gnd DFFSR_175/S FILL
XINVX1_201 BUFX2_73/A OR2X2_6/gnd INVX1_201/Y DFFSR_92/S INVX1
XFILL_8_NAND3X1_194 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_7_NAND3X1_24 INVX1_1/gnd DFFSR_97/S FILL
XFILL_1_DFFSR_224 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_4_BUFX2_34 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_28_DFFSR_151 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_4_DFFPOSX1_13 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_42_DFFSR_255 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_1_NAND2X1_175 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_6_NAND3X1_27 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_18_DFFSR_154 BUFX2_99/A DFFSR_7/S FILL
XFILL_32_DFFSR_258 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_6_OAI22X1_12 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_5_NAND3X1_30 BUFX2_79/A DFFSR_6/S FILL
XNAND3X1_27 BUFX2_85/A AND2X2_3/Y BUFX2_21/Y OR2X2_4/gnd AND2X2_9/A DFFSR_3/S NAND3X1
XFILL_53_4_0 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_22_DFFSR_261 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_5_OAI22X1_15 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_4_NAND3X1_33 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_41_DFFSR_56 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_30_DFFSR_96 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_2_INVX1_90 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_3_NOR2X1_33 INVX1_3/gnd DFFSR_23/S FILL
XFILL_13_DFFPOSX1_32 INVX1_67/gnd DFFSR_201/S FILL
XOAI22X1_12 INVX1_28/Y OAI22X1_6/B INVX1_29/Y OAI22X1_6/D DFFSR_28/gnd NOR2X1_16/A
+ DFFSR_3/S OAI22X1
XFILL_12_DFFSR_264 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_4_OAI22X1_18 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_3_NAND3X1_36 DFFSR_8/gnd DFFSR_8/S FILL
XDFFSR_154 INVX1_74/A CLKBUF1_3/Y BUFX2_63/Y DFFSR_7/S DFFSR_154/D BUFX2_99/A DFFSR_7/S
+ DFFSR
XFILL_2_NAND2X1_109 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_51_6_1 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_2_NAND3X1_39 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_3_OAI22X1_21 BUFX2_98/A DFFSR_32/S FILL
XFILL_8_DFFSR_13 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_4_DFFSR_151 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_14_DFFSR_46 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_2_OAI22X1_24 BUFX2_98/A DFFSR_32/S FILL
XFILL_1_NAND3X1_42 BUFX2_79/A DFFSR_6/S FILL
XFILL_1_BUFX2_81 BUFX2_79/A DFFSR_7/S FILL
XFILL_45_DFFSR_182 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_1_OAI22X1_27 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_0_NAND3X1_45 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_8_DFFSR_258 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_35_DFFSR_185 INVX1_39/gnd DFFSR_54/S FILL
XFILL_23_DFFPOSX1_21 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_0_OAI22X1_30 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_25_DFFSR_188 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_49_DFFSR_63 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_15_DFFSR_191 INVX1_67/gnd DFFSR_175/S FILL
XFILL_7_NAND3X1_224 INVX1_39/gnd DFFSR_54/S FILL
XFILL_3_DFFPOSX1_43 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_5_DFFSR_60 OR2X2_3/gnd DFFSR_60/S FILL
XINVX1_47 INVX1_47/A BUFX2_77/gnd INVX1_47/Y DFFSR_98/S INVX1
XFILL_11_DFFSR_93 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_33_DFFSR_13 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_22_DFFSR_53 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_0_NOR2X1_70 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_48_DFFSR_109 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_38_DFFSR_112 OR2X2_4/gnd DFFSR_32/S FILL
XINVX1_165 BUFX2_99/A BUFX2_99/A NOR2X1_69/B DFFSR_92/S INVX1
XFILL_8_NAND3X1_158 AND2X2_38/B DFFSR_59/S FILL
XFILL_1_DFFSR_188 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_28_DFFSR_115 INVX1_1/gnd DFFSR_97/S FILL
XFILL_42_DFFSR_219 INVX1_67/gnd DFFSR_175/S FILL
XFILL_1_NAND2X1_139 INVX1_1/gnd DFFSR_97/S FILL
XFILL_4_INVX1_162 INVX1_39/gnd DFFSR_34/S FILL
XFILL_7_AND2X2_29 AND2X2_38/B DFFSR_23/S FILL
XFILL_18_DFFSR_118 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_32_DFFSR_222 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_1_NAND2X1_9 BUFX2_79/A DFFSR_6/S FILL
XFILL_22_DFFSR_225 INVX1_67/gnd DFFSR_175/S FILL
XFILL_30_DFFSR_60 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_2_INVX1_54 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_41_DFFSR_20 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_12_DFFSR_228 XOR2X1_1/gnd DFFSR_208/S FILL
XDFFSR_118 INVX1_44/A DFFSR_57/CLK DFFSR_35/R DFFSR_60/S DFFSR_118/D OR2X2_3/gnd DFFSR_60/S
+ DFFSR
XFILL_14_DFFSR_10 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_4_DFFSR_115 INVX1_1/gnd DFFSR_97/S FILL
XFILL_1_BUFX2_45 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_1_OAI22X1_8 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_45_DFFSR_146 BUFX2_79/A DFFSR_7/S FILL
XFILL_8_DFFSR_222 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_8_DFFSR_3 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_35_DFFSR_149 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_49_DFFSR_253 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_25_DFFSR_152 INVX1_1/gnd DFFSR_53/S FILL
XFILL_49_DFFSR_27 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_39_DFFSR_256 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_1_INVX1_199 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_38_DFFSR_67 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_15_DFFSR_155 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_7_NAND3X1_188 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_29_DFFSR_259 BUFX2_79/A DFFSR_6/S FILL
XINVX1_11 DFFSR_58/Q OR2X2_3/gnd INVX1_11/Y DFFSR_4/S INVX1
XFILL_0_NAND2X1_169 INVX1_1/gnd DFFSR_53/S FILL
XDFFSR_64 DFFSR_56/D CLKBUF1_37/Y DFFSR_8/R DFFSR_60/S DFFSR_48/Q OR2X2_3/gnd DFFSR_60/S
+ DFFSR
XFILL_19_DFFSR_262 BUFX2_98/A DFFSR_32/S FILL
XFILL_5_DFFSR_24 BUFX2_98/A DFFSR_6/S FILL
XFILL_22_DFFSR_17 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_11_DFFSR_57 BUFX2_79/A DFFSR_6/S FILL
XFILL_0_NOR2X1_34 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_27_2_0 INVX1_3/gnd DFFSR_79/S FILL
XFILL_6_OR2X2_3 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_8_NAND3X1_122 XOR2X1_4/gnd DFFSR_97/S FILL
XINVX1_129 BUFX2_35/Y AND2X2_38/B INVX1_129/Y DFFSR_23/S INVX1
XFILL_4_NOR2X1_5 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_1_DFFSR_152 INVX1_1/gnd DFFSR_53/S FILL
XFILL_12_DFFPOSX1_26 AND2X2_38/B DFFSR_23/S FILL
XFILL_25_4_1 AND2X2_38/B DFFSR_23/S FILL
XFILL_32_DFFSR_7 BUFX2_79/A DFFSR_7/S FILL
XFILL_1_NAND2X1_103 AND2X2_38/B DFFSR_23/S FILL
XFILL_42_DFFSR_183 INVX1_67/gnd DFFSR_175/S FILL
XFILL_46_DFFSR_74 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_7_3_0 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_5_DFFSR_259 BUFX2_79/A DFFSR_6/S FILL
XFILL_32_DFFSR_186 BUFX2_99/A DFFSR_92/S FILL
XFILL_23_6_2 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_22_DFFSR_189 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_30_DFFSR_24 BUFX2_98/A DFFSR_6/S FILL
XFILL_2_DFFSR_71 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_2_INVX1_18 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_5_5_1 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_19_DFFSR_64 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_6_BUFX2_99 BUFX2_99/A DFFSR_7/S FILL
XFILL_12_DFFSR_192 INVX1_1/gnd DFFSR_97/S FILL
XFILL_22_DFFPOSX1_15 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_6_NAND3X1_218 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_6_XOR2X1_1 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_45_DFFSR_110 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_2_DFFPOSX1_37 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_8_DFFSR_186 BUFX2_99/A DFFSR_92/S FILL
XFILL_35_DFFSR_113 BUFX2_99/A DFFSR_92/S FILL
XAND2X2_33 INVX1_135/A AND2X2_33/B NOR3X1_6/gnd AND2X2_33/Y DFFSR_79/S AND2X2
XFILL_49_DFFSR_217 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_25_DFFSR_116 INVX1_3/gnd DFFSR_23/S FILL
XFILL_39_DFFSR_220 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_1_INVX1_163 INVX1_39/gnd DFFSR_54/S FILL
XFILL_4_AND2X2_30 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_38_DFFSR_31 BUFX2_79/A DFFSR_6/S FILL
XFILL_27_DFFSR_71 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_15_DFFSR_119 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_7_NAND3X1_152 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_29_DFFSR_223 INVX1_39/gnd DFFSR_34/S FILL
XFILL_0_NAND2X1_133 BUFX2_72/gnd DFFSR_201/S FILL
XDFFSR_28 DFFSR_28/Q DFFSR_8/CLK DFFSR_2/R DFFSR_8/S DFFSR_4/Q DFFSR_28/gnd DFFSR_8/S
+ DFFSR
XFILL_19_DFFSR_226 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_11_DFFSR_21 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_8_OAI22X1_6 BUFX2_98/A DFFSR_32/S FILL
XFILL_2_NOR3X1_2 INVX1_1/gnd DFFSR_53/S FILL
XFILL_1_DFFSR_116 INVX1_3/gnd DFFSR_23/S FILL
XFILL_17_5 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_33_1_2 INVX1_1/gnd DFFSR_53/S FILL
XFILL_21_DFFPOSX1_45 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_42_DFFSR_147 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_35_DFFSR_78 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_46_DFFSR_38 BUFX2_98/A DFFSR_6/S FILL
XFILL_5_DFFSR_223 INVX1_39/gnd DFFSR_34/S FILL
XFILL_32_DFFSR_150 AND2X2_38/B DFFSR_23/S FILL
XFILL_5_NAND3X1_248 INVX1_3/gnd DFFSR_79/S FILL
XFILL_46_DFFSR_254 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_22_DFFSR_153 INVX1_67/gnd DFFSR_201/S FILL
XFILL_2_DFFSR_35 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_36_DFFSR_257 INVX1_39/gnd DFFSR_34/S FILL
XFILL_19_DFFSR_28 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_12_DFFSR_156 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_6_BUFX2_63 BUFX2_98/A DFFSR_32/S FILL
XFILL_26_DFFSR_260 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_8_OAI21X1_104 INVX1_67/gnd DFFSR_201/S FILL
XFILL_16_DFFSR_263 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_20_CLKBUF1_18 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_6_NAND3X1_182 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_19_CLKBUF1_21 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_19_DFFSR_1 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_43_DFFSR_85 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_8_DFFSR_150 AND2X2_38/B DFFSR_23/S FILL
XFILL_18_CLKBUF1_24 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_49_DFFSR_181 INVX1_3/gnd DFFSR_79/S FILL
XNAND3X1_218 NAND3X1_187/Y NAND3X1_218/B XOR2X1_8/A DFFSR_46/gnd NAND3X1_218/Y DFFSR_54/S
+ NAND3X1
XFILL_17_CLKBUF1_27 INVX1_1/gnd DFFSR_97/S FILL
XFILL_39_DFFSR_184 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_1_INVX1_127 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_27_DFFSR_35 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_16_DFFSR_75 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_2_DFFSR_260 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_7_NAND3X1_116 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_16_CLKBUF1_30 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_29_DFFSR_187 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_3_BUFX2_2 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_11_DFFPOSX1_20 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_19_DFFSR_190 INVX1_39/gnd DFFSR_34/S FILL
XFILL_15_CLKBUF1_33 XOR2X1_4/gnd DFFSR_91/S FILL
XNOR2X1_72 INVX1_175/Y INVX1_161/Y DFFSR_8/gnd NOR2X1_72/Y DFFSR_60/S NOR2X1
XFILL_14_CLKBUF1_36 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_51_DFFSR_92 BUFX2_99/A DFFSR_92/S FILL
XFILL_4_NOR2X1_69 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_13_CLKBUF1_39 INVX1_1/gnd DFFSR_53/S FILL
XFILL_12_CLKBUF1_42 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_42_DFFSR_111 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_35_DFFSR_42 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_7_DFFSR_89 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_24_DFFSR_82 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_11_CLKBUF1_45 BUFX2_79/A DFFSR_7/S FILL
XFILL_5_DFFSR_187 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_32_DFFSR_114 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_46_DFFSR_218 BUFX2_98/A DFFSR_32/S FILL
XFILL_10_CLKBUF1_48 INVX1_3/gnd DFFSR_79/S FILL
XFILL_5_NAND3X1_212 INVX1_39/gnd DFFSR_54/S FILL
XFILL_22_DFFSR_117 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_1_DFFPOSX1_31 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_36_DFFSR_221 AND2X2_38/B DFFSR_59/S FILL
XFILL_1_AND2X2_31 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_12_DFFSR_120 INVX1_3/gnd DFFSR_23/S FILL
XFILL_5_NAND2X1_8 INVX1_1/gnd DFFSR_53/S FILL
XFILL_6_BUFX2_27 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_26_DFFSR_224 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_16_DFFSR_227 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_16_NOR3X1_6 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_6_NAND3X1_146 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_10_DFFPOSX1_50 INVX1_1/gnd DFFSR_53/S FILL
XFILL_43_DFFSR_49 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_8_DFFSR_114 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_32_DFFSR_89 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_5_OAI22X1_7 AND2X2_38/B DFFSR_59/S FILL
XFILL_49_DFFSR_145 BUFX2_72/gnd DFFSR_201/S FILL
XNAND3X1_182 INVX1_158/Y OAI21X1_48/Y OAI21X1_49/Y DFFSR_34/gnd AOI22X1_24/B DFFSR_1/S
+ NAND3X1
XFILL_39_DFFSR_148 INVX1_67/gnd DFFSR_175/S FILL
XFILL_16_DFFSR_39 INVX1_3/gnd DFFSR_79/S FILL
XFILL_3_BUFX2_74 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_2_DFFSR_224 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_29_DFFSR_151 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_43_DFFSR_255 OR2X2_4/gnd DFFSR_32/S FILL
XNAND3X1_1 DFFSR_57/D BUFX2_16/Y BUFX2_14/Y BUFX2_98/A NAND3X1_4/B DFFSR_6/S NAND3X1
XFILL_20_DFFPOSX1_39 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_19_DFFSR_154 BUFX2_99/A DFFSR_7/S FILL
XFILL_33_DFFSR_258 DFFSR_5/gnd DFFSR_5/S FILL
XNOR2X1_36 NOR3X1_4/A NOR3X1_4/B OR2X2_1/gnd BUFX2_27/A DFFSR_51/S NOR2X1
XFILL_4_NAND3X1_242 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_23_DFFSR_261 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_40_DFFSR_96 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_4_NOR2X1_33 INVX1_3/gnd DFFSR_23/S FILL
XFILL_13_DFFSR_264 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_1_AND2X2_5 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_7_DFFSR_53 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_5_DFFSR_151 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_13_DFFSR_86 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_24_DFFSR_46 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_5_NAND3X1_176 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_10_CLKBUF1_12 AND2X2_38/B DFFSR_23/S FILL
XFILL_46_DFFSR_182 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_9_DFFSR_258 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_36_DFFSR_185 INVX1_39/gnd DFFSR_54/S FILL
XFILL_26_DFFSR_188 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_34_2_0 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_9_CLKBUF1_15 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_16_DFFSR_191 INVX1_67/gnd DFFSR_175/S FILL
XFILL_10_DFFSR_8 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_8_CLKBUF1_18 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_6_NAND3X1_110 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_7_CLKBUF1_21 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_32_4_1 INVX1_1/gnd DFFSR_97/S FILL
XFILL_10_DFFPOSX1_14 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_21_DFFSR_93 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_43_DFFSR_13 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_32_DFFSR_53 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_1_NOR2X1_70 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_6_CLKBUF1_24 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_49_DFFSR_109 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_5_CLKBUF1_27 INVX1_1/gnd DFFSR_97/S FILL
XNAND3X1_146 INVX1_144/A AOI22X1_19/C OAI21X1_38/C BUFX2_8/gnd AOI21X1_14/A DFFSR_51/S
+ NAND3X1
XFILL_30_6_2 XOR2X1_4/gnd DFFSR_91/S FILL
XCLKBUF1_24 BUFX2_2/Y DFFSR_4/gnd DFFSR_93/CLK DFFSR_98/S CLKBUF1
XFILL_39_DFFSR_112 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_4_CLKBUF1_30 BUFX2_77/gnd DFFSR_5/S FILL
XOR2X2_4 OR2X2_4/A OR2X2_4/B OR2X2_4/gnd OR2X2_4/Y DFFSR_32/S OR2X2
XFILL_3_BUFX2_38 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_2_DFFSR_188 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_29_DFFSR_115 INVX1_1/gnd DFFSR_97/S FILL
XFILL_43_DFFSR_219 INVX1_67/gnd DFFSR_175/S FILL
XFILL_3_CLKBUF1_33 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_8_AND2X2_29 AND2X2_38/B DFFSR_23/S FILL
XFILL_19_DFFSR_118 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_33_DFFSR_222 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_2_CLKBUF1_36 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_31_DFFSR_4 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_2_NAND2X1_9 BUFX2_79/A DFFSR_6/S FILL
XFILL_23_DFFSR_225 INVX1_67/gnd DFFSR_175/S FILL
XFILL_1_CLKBUF1_39 INVX1_1/gnd DFFSR_53/S FILL
XFILL_4_NAND3X1_206 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_1_INVX1_94 INVX1_67/gnd DFFSR_201/S FILL
XFILL_40_DFFSR_60 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_0_CLKBUF1_42 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_0_DFFPOSX1_25 BUFX2_79/A DFFSR_6/S FILL
XFILL_13_DFFSR_228 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_7_DFFSR_17 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_24_DFFSR_10 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_13_DFFSR_50 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_5_DFFSR_115 INVX1_1/gnd DFFSR_97/S FILL
XFILL_0_BUFX2_85 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_2_OAI22X1_8 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_46_DFFSR_146 BUFX2_79/A DFFSR_7/S FILL
XFILL_5_NAND3X1_140 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_9_DFFSR_222 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_36_DFFSR_149 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_50_DFFSR_253 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_26_DFFSR_152 INVX1_1/gnd DFFSR_53/S FILL
XFILL_40_DFFSR_256 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_48_DFFSR_67 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_2_INVX1_199 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_16_DFFSR_155 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_30_DFFSR_259 BUFX2_79/A DFFSR_6/S FILL
XFILL_20_DFFSR_262 BUFX2_98/A DFFSR_32/S FILL
XFILL_32_DFFSR_17 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_4_DFFSR_64 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_4_INVX1_11 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_21_DFFSR_57 BUFX2_79/A DFFSR_6/S FILL
XFILL_40_1_2 BUFX2_98/A DFFSR_6/S FILL
XFILL_10_DFFSR_97 INVX1_1/gnd DFFSR_97/S FILL
XFILL_19_DFFPOSX1_33 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_1_NOR2X1_34 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_10_DFFSR_265 INVX1_67/gnd DFFSR_175/S FILL
XNAND3X1_110 DFFSR_206/D BUFX2_27/Y NOR2X1_31/Y XOR2X1_1/gnd NAND3X1_110/Y DFFSR_151/S
+ NAND3X1
XFILL_3_NAND3X1_236 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_2_DFFSR_152 INVX1_1/gnd DFFSR_53/S FILL
XFILL_43_DFFSR_183 INVX1_67/gnd DFFSR_175/S FILL
XFILL_6_DFFSR_259 BUFX2_79/A DFFSR_6/S FILL
XFILL_33_DFFSR_186 BUFX2_99/A DFFSR_92/S FILL
XFILL_23_DFFSR_189 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_4_NAND3X1_170 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_40_DFFSR_24 BUFX2_98/A DFFSR_6/S FILL
XFILL_1_INVX1_58 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_29_DFFSR_64 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_13_DFFSR_192 INVX1_1/gnd DFFSR_97/S FILL
XFILL_9_DFFPOSX1_44 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_13_DFFSR_14 INVX1_1/gnd DFFSR_53/S FILL
XFILL_0_BUFX2_49 INVX1_1/gnd DFFSR_97/S FILL
XFILL_46_DFFSR_110 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_5_NAND3X1_104 AND2X2_38/B DFFSR_23/S FILL
XFILL_9_DFFSR_186 BUFX2_99/A DFFSR_92/S FILL
XFILL_36_DFFSR_113 BUFX2_99/A DFFSR_92/S FILL
XFILL_50_DFFSR_217 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_26_DFFSR_116 INVX1_3/gnd DFFSR_23/S FILL
XFILL_40_DFFSR_220 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_48_DFFSR_31 BUFX2_79/A DFFSR_6/S FILL
XFILL_37_DFFSR_71 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_2_INVX1_163 INVX1_39/gnd DFFSR_54/S FILL
XFILL_5_AND2X2_30 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_16_DFFSR_119 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_30_DFFSR_223 INVX1_39/gnd DFFSR_34/S FILL
XFILL_20_DFFSR_226 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_4_DFFSR_28 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_21_DFFSR_21 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_10_DFFSR_61 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_10_DFFSR_229 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_3_NAND3X1_200 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_9_OAI22X1_6 BUFX2_98/A DFFSR_32/S FILL
XFILL_3_NOR2X1_9 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_2_DFFSR_116 INVX1_3/gnd DFFSR_23/S FILL
XFILL_43_DFFSR_147 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_45_DFFSR_78 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_6_DFFSR_223 INVX1_39/gnd DFFSR_34/S FILL
XFILL_33_DFFSR_150 AND2X2_38/B DFFSR_23/S FILL
XFILL_47_DFFSR_254 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_23_DFFSR_153 INVX1_67/gnd DFFSR_201/S FILL
XFILL_4_NAND3X1_134 INVX1_39/gnd DFFSR_54/S FILL
XFILL_1_INVX1_22 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_1_DFFSR_75 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_37_DFFSR_257 INVX1_39/gnd DFFSR_34/S FILL
XFILL_29_DFFSR_28 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_18_DFFSR_68 BUFX2_98/A DFFSR_6/S FILL
XFILL_13_DFFSR_156 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_27_DFFSR_260 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_6_NAND2X1_170 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_17_DFFSR_263 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_0_BUFX2_13 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_5_XOR2X1_5 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_21_DFFPOSX1_3 INVX1_39/gnd DFFSR_34/S FILL
XFILL_9_DFFSR_150 AND2X2_38/B DFFSR_23/S FILL
XFILL_43_DFFSR_7 BUFX2_79/A DFFSR_7/S FILL
XFILL_20_DFFPOSX1_6 AND2X2_38/B DFFSR_23/S FILL
XFILL_18_DFFPOSX1_27 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_50_DFFSR_181 INVX1_3/gnd DFFSR_79/S FILL
XFILL_19_DFFPOSX1_9 INVX1_67/gnd DFFSR_201/S FILL
XFILL_40_DFFSR_184 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_2_INVX1_127 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_37_DFFSR_35 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_9_DFFSR_82 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_26_DFFSR_75 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_2_NAND3X1_230 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_3_DFFSR_260 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_30_DFFSR_187 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_20_DFFSR_190 INVX1_39/gnd DFFSR_34/S FILL
XFILL_10_DFFSR_25 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_10_DFFSR_193 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_5_NOR2X1_69 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_3_NAND3X1_164 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_1_NOR3X1_6 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_43_DFFSR_111 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_8_DFFPOSX1_38 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_34_DFFSR_82 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_45_DFFSR_42 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_41_2_0 BUFX2_98/A DFFSR_32/S FILL
XFILL_6_DFFSR_187 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_33_DFFSR_114 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_47_DFFSR_218 BUFX2_98/A DFFSR_32/S FILL
XFILL_23_DFFSR_117 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_1_DFFSR_39 INVX1_3/gnd DFFSR_79/S FILL
XFILL_37_DFFSR_221 AND2X2_38/B DFFSR_59/S FILL
XFILL_18_DFFSR_32 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_39_4_1 BUFX2_79/A DFFSR_6/S FILL
XFILL_2_AND2X2_31 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_5_BUFX2_67 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_6_NAND2X1_8 INVX1_1/gnd DFFSR_53/S FILL
XFILL_13_DFFSR_120 INVX1_3/gnd DFFSR_23/S FILL
XFILL_27_DFFSR_224 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_6_NAND2X1_134 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_17_DFFSR_227 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_37_6_2 BUFX2_99/A DFFSR_7/S FILL
XXOR2X1_9 XOR2X1_9/A XOR2X1_9/B NOR3X1_6/gnd XOR2X1_9/Y DFFSR_79/S XOR2X1
XFILL_11_XOR2X1_2 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_9_DFFSR_114 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_42_DFFSR_89 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_9_AOI21X1_59 OR2X2_1/gnd DFFSR_51/S FILL
XNAND2X1_170 DFFSR_216/S DFFPOSX1_37/Q BUFX2_7/gnd NOR2X1_74/B DFFSR_216/S NAND2X1
XFILL_6_OAI22X1_7 AND2X2_38/B DFFSR_59/S FILL
XFILL_50_DFFSR_145 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_4_OAI21X1_116 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_8_AOI21X1_62 INVX1_3/gnd DFFSR_23/S FILL
XFILL_27_DFFPOSX1_46 INVX1_39/gnd DFFSR_34/S FILL
XFILL_40_DFFSR_148 INVX1_67/gnd DFFSR_175/S FILL
XFILL_26_DFFSR_39 INVX1_3/gnd DFFSR_79/S FILL
XFILL_7_AOI21X1_65 INVX1_3/gnd DFFSR_23/S FILL
XFILL_9_DFFSR_46 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_15_DFFSR_79 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_2_NAND3X1_194 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_3_DFFSR_224 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_30_DFFSR_151 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_6_AOI21X1_68 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_44_DFFSR_255 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_20_DFFSR_154 BUFX2_99/A DFFSR_7/S FILL
XFILL_34_DFFSR_258 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_5_AOI21X1_71 BUFX2_99/A DFFSR_92/S FILL
XAOI21X1_68 AOI21X1_68/A AOI21X1_66/Y AOI21X1_68/C XOR2X1_4/gnd OR2X2_6/A DFFSR_97/S
+ AOI21X1
XFILL_10_DFFSR_157 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_24_DFFSR_261 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_50_DFFSR_96 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_3_NAND3X1_128 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_5_NOR2X1_33 INVX1_3/gnd DFFSR_23/S FILL
XFILL_30_DFFSR_1 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_14_DFFSR_264 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_5_NAND2X1_164 INVX1_67/gnd DFFSR_175/S FILL
XFILL_6_DFFSR_93 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_23_DFFSR_86 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_34_DFFSR_46 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_6_DFFSR_151 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_47_DFFSR_182 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_37_DFFSR_185 INVX1_39/gnd DFFSR_54/S FILL
XBUFX2_71 BUFX2_71/A DFFSR_5/gnd dout[0] DFFSR_5/S BUFX2
XFILL_0_DFFSR_261 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_5_BUFX2_31 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_17_DFFPOSX1_21 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_47_1_2 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_27_DFFSR_188 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_17_DFFSR_191 INVX1_67/gnd DFFSR_175/S FILL
XFILL_1_NAND3X1_224 INVX1_39/gnd DFFSR_54/S FILL
XFILL_9_DFFPOSX1_3 INVX1_39/gnd DFFSR_34/S FILL
XFILL_3_INVX1_87 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_42_DFFSR_53 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_8_DFFPOSX1_6 AND2X2_38/B DFFSR_23/S FILL
XFILL_31_DFFSR_93 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_9_AOI21X1_23 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_2_NOR2X1_70 XOR2X1_4/gnd DFFSR_91/S FILL
XNAND2X1_134 DFFSR_1/S INVX1_192/A DFFSR_1/gnd NAND2X1_134/Y DFFSR_1/S NAND2X1
XFILL_50_DFFSR_109 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_7_DFFPOSX1_9 INVX1_67/gnd DFFSR_201/S FILL
XFILL_27_DFFPOSX1_10 INVX1_67/gnd DFFSR_201/S FILL
XFILL_8_AOI21X1_26 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_40_DFFSR_112 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_9_DFFSR_10 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_7_AOI21X1_29 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_15_DFFSR_43 BUFX2_98/A DFFSR_6/S FILL
XFILL_2_NAND3X1_158 AND2X2_38/B DFFSR_59/S FILL
XFILL_3_DFFSR_188 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_2_BUFX2_78 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_30_DFFSR_115 INVX1_1/gnd DFFSR_97/S FILL
XFILL_15_0_0 INVX1_39/gnd DFFSR_34/S FILL
XFILL_6_AOI21X1_32 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_44_DFFSR_219 INVX1_67/gnd DFFSR_175/S FILL
XFILL_7_DFFPOSX1_32 INVX1_67/gnd DFFSR_201/S FILL
XFILL_20_DFFSR_118 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_34_DFFSR_222 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_5_AOI21X1_35 INVX1_39/gnd DFFSR_54/S FILL
XAOI21X1_32 AOI21X1_32/A AOI21X1_32/B OAI21X1_53/C DFFSR_62/gnd AOI21X1_33/C DFFSR_208/S
+ AOI21X1
XFILL_3_NAND2X1_9 BUFX2_79/A DFFSR_6/S FILL
XFILL_10_DFFSR_121 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_4_AOI21X1_38 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_13_2_1 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_24_DFFSR_225 INVX1_67/gnd DFFSR_175/S FILL
XFILL_50_DFFSR_60 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_3_AOI21X1_41 INVX1_39/gnd DFFSR_34/S FILL
XFILL_14_DFFSR_228 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_2_AOI21X1_44 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_11_4_2 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_0_AND2X2_9 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_5_NAND2X1_128 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_34_DFFSR_10 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_23_DFFSR_50 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_12_DFFSR_90 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_6_DFFSR_57 BUFX2_79/A DFFSR_6/S FILL
XFILL_1_AOI21X1_47 INVX1_67/gnd DFFSR_175/S FILL
XFILL_6_DFFSR_115 INVX1_1/gnd DFFSR_97/S FILL
XFILL_3_OAI22X1_8 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_47_DFFSR_146 BUFX2_79/A DFFSR_7/S FILL
XFILL_0_AOI21X1_50 INVX1_67/gnd DFFSR_175/S FILL
XFILL_37_DFFSR_149 BUFX2_72/gnd DFFSR_276/S FILL
XBUFX2_35 rst OR2X2_1/gnd BUFX2_35/Y DFFSR_59/S BUFX2
XFILL_0_DFFSR_225 INVX1_67/gnd DFFSR_175/S FILL
XFILL_27_DFFSR_152 INVX1_1/gnd DFFSR_53/S FILL
XFILL_3_OAI21X1_110 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_41_DFFSR_256 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_9_OAI21X1_71 INVX1_3/gnd DFFSR_79/S FILL
XFILL_26_DFFPOSX1_40 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_3_INVX1_199 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_17_DFFSR_155 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_8_OAI21X1_74 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_1_NAND3X1_188 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_31_DFFSR_259 BUFX2_79/A DFFSR_6/S FILL
XFILL_7_OAI21X1_77 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_6_NAND2X1_95 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_21_DFFSR_262 BUFX2_98/A DFFSR_32/S FILL
XFILL_42_DFFSR_17 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_3_INVX1_51 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_31_DFFSR_57 BUFX2_79/A DFFSR_6/S FILL
XFILL_20_DFFSR_97 INVX1_1/gnd DFFSR_97/S FILL
XFILL_2_NOR2X1_34 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_11_DFFSR_265 INVX1_67/gnd DFFSR_175/S FILL
XFILL_6_OAI21X1_80 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_5_NAND2X1_98 OR2X2_6/gnd DFFSR_53/S FILL
XNAND2X1_95 AND2X2_34/B AND2X2_35/B XOR2X1_4/gnd XNOR2X1_3/A DFFSR_91/S NAND2X1
XFILL_5_OAI21X1_83 DFFSR_34/gnd DFFSR_1/S FILL
XOAI21X1_80 OAI21X1_80/A OAI21X1_80/B INVX1_179/A OR2X2_3/gnd AOI21X1_38/B DFFSR_60/S
+ OAI21X1
XFILL_2_NAND3X1_122 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_4_OAI21X1_86 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_3_DFFSR_152 INVX1_1/gnd DFFSR_53/S FILL
XFILL_2_BUFX2_42 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_44_DFFSR_183 INVX1_67/gnd DFFSR_175/S FILL
XFILL_3_OAI21X1_89 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_7_DFFSR_259 BUFX2_79/A DFFSR_6/S FILL
XFILL_34_DFFSR_186 BUFX2_99/A DFFSR_92/S FILL
XFILL_4_NAND2X1_158 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_21_DFFSR_8 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_2_OAI21X1_92 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_24_DFFSR_189 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_1_OAI21X1_95 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_39_DFFSR_64 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_50_DFFSR_24 BUFX2_98/A DFFSR_6/S FILL
XFILL_0_INVX1_98 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_14_DFFSR_192 INVX1_1/gnd DFFSR_97/S FILL
XFILL_0_OAI21X1_98 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_16_DFFPOSX1_15 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_6_DFFSR_21 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_23_DFFSR_14 INVX1_1/gnd DFFSR_53/S FILL
XFILL_12_DFFSR_54 INVX1_39/gnd DFFSR_54/S FILL
XFILL_5_BUFX2_9 AND2X2_38/B DFFSR_59/S FILL
XFILL_1_AOI21X1_11 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_47_DFFSR_110 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_0_NAND3X1_218 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_1_0_2 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_0_AOI21X1_14 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_37_DFFSR_113 BUFX2_99/A DFFSR_92/S FILL
XFILL_51_DFFSR_217 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_5_NOR2X1_2 INVX1_1/gnd DFFSR_97/S FILL
XFILL_0_DFFSR_189 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_27_DFFSR_116 INVX1_3/gnd DFFSR_23/S FILL
XFILL_42_DFFSR_4 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_41_DFFSR_220 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_47_DFFSR_71 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_3_INVX1_163 INVX1_39/gnd DFFSR_54/S FILL
XFILL_6_AND2X2_30 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_17_DFFSR_119 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_8_OAI21X1_38 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_1_NAND3X1_152 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_31_DFFSR_223 INVX1_39/gnd DFFSR_34/S FILL
XFILL_7_OAI21X1_41 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_6_NAND2X1_59 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_21_DFFSR_226 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_31_DFFSR_21 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_3_INVX1_15 BUFX2_98/A DFFSR_32/S FILL
XFILL_3_DFFSR_68 BUFX2_98/A DFFSR_6/S FILL
XFILL_20_DFFSR_61 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_6_DFFPOSX1_26 AND2X2_38/B DFFSR_23/S FILL
XFILL_5_NAND2X1_62 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_48_2_0 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_11_DFFSR_229 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_6_OAI21X1_44 DFFSR_62/gnd DFFSR_208/S FILL
XNAND2X1_59 NAND2X1_59/A INVX1_131/Y DFFSR_62/gnd XOR2X1_1/A DFFSR_208/S NAND2X1
XFILL_4_NAND2X1_65 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_5_OAI21X1_47 DFFSR_34/gnd DFFSR_1/S FILL
XOAI21X1_44 AOI21X1_19/Y INVX1_156/Y AOI21X1_18/Y DFFSR_62/gnd OAI21X1_44/Y DFFSR_208/S
+ OAI21X1
XFILL_4_OAI21X1_50 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_3_DFFSR_116 INVX1_3/gnd DFFSR_23/S FILL
XFILL_3_NAND2X1_68 AND2X2_38/B DFFSR_23/S FILL
XFILL_46_4_1 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_0_OAI22X1_9 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_44_DFFSR_147 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_15_DFFPOSX1_45 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_2_NAND2X1_71 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_3_OAI21X1_53 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_7_DFFSR_223 INVX1_39/gnd DFFSR_34/S FILL
XFILL_4_NAND2X1_122 INVX1_67/gnd DFFSR_175/S FILL
XFILL_34_DFFSR_150 AND2X2_38/B DFFSR_23/S FILL
XFILL_1_NAND2X1_74 AND2X2_38/B DFFSR_59/S FILL
XFILL_48_DFFSR_254 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_2_OAI21X1_56 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_44_6_2 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_11_AOI22X1_22 INVX1_3/gnd DFFSR_79/S FILL
XFILL_24_DFFSR_153 INVX1_67/gnd DFFSR_201/S FILL
XFILL_0_NAND2X1_77 AND2X2_38/B DFFSR_23/S FILL
XFILL_38_DFFSR_257 INVX1_39/gnd DFFSR_34/S FILL
XFILL_1_OAI21X1_59 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_0_INVX1_200 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_39_DFFSR_28 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_28_DFFSR_68 BUFX2_98/A DFFSR_6/S FILL
XFILL_10_AOI22X1_25 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_0_INVX1_62 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_14_DFFSR_156 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_0_OAI21X1_62 INVX1_3/gnd DFFSR_79/S FILL
XFILL_28_DFFSR_260 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_2_OAI21X1_104 INVX1_67/gnd DFFSR_201/S FILL
XFILL_25_DFFPOSX1_34 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_18_DFFSR_263 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_9_AOI22X1_28 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_12_DFFSR_18 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_0_NAND3X1_182 DFFSR_34/gnd DFFSR_1/S FILL
XNOR2X1_6 NOR2X1_6/A NOR2X1_6/B BUFX2_98/A NOR2X1_6/Y DFFSR_6/S NOR2X1
XFILL_0_DFFSR_153 INVX1_67/gnd DFFSR_201/S FILL
XDFFSR_263 DFFSR_7/D CLKBUF1_8/Y DFFSR_257/R DFFSR_51/S DFFSR_263/D OR2X2_1/gnd DFFSR_51/S
+ DFFSR
XFILL_12_5_0 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_41_DFFSR_184 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_47_DFFSR_35 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_3_INVX1_127 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_36_DFFSR_75 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_4_DFFSR_260 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_31_DFFSR_187 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_1_NAND3X1_116 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_6_NAND2X1_23 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_21_DFFSR_190 INVX1_39/gnd DFFSR_34/S FILL
XFILL_3_DFFSR_32 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_20_DFFSR_25 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_5_NAND2X1_26 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_11_DFFSR_193 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_3_NAND2X1_152 INVX1_1/gnd DFFSR_97/S FILL
XNAND2X1_23 DFFSR_119/D NOR2X1_5/Y DFFSR_8/gnd OAI21X1_7/C DFFSR_8/S NAND2X1
XFILL_4_NAND2X1_29 INVX1_3/gnd DFFSR_23/S FILL
XFILL_5_OAI21X1_11 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_6_NOR2X1_69 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_8_3 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_3_NAND2X1_32 INVX1_3/gnd DFFSR_79/S FILL
XFILL_4_OAI21X1_14 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_9_DFFSR_7 BUFX2_79/A DFFSR_7/S FILL
XDFFPOSX1_26 NAND2X1_156/A CLKBUF1_45/Y AOI21X1_54/Y AND2X2_38/B DFFSR_23/S DFFPOSX1
XFILL_44_DFFSR_111 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_2_NAND2X1_35 INVX1_67/gnd DFFSR_201/S FILL
XFILL_54_1_2 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_3_OAI21X1_17 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_44_DFFSR_82 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_7_DFFSR_187 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_34_DFFSR_114 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_9_NAND3X1_91 AND2X2_38/B DFFSR_59/S FILL
XFILL_48_DFFSR_218 BUFX2_98/A DFFSR_32/S FILL
XFILL_2_OAI21X1_20 AND2X2_38/B DFFSR_23/S FILL
XFILL_1_NAND2X1_38 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_24_DFFSR_117 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_8_NAND3X1_94 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_1_OAI21X1_23 INVX1_67/gnd DFFSR_201/S FILL
XFILL_0_NAND2X1_41 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_38_DFFSR_221 AND2X2_38/B DFFSR_59/S FILL
XAOI21X1_2 AOI21X1_2/A INVX1_120/Y BUFX2_39/Y DFFSR_62/gnd AOI21X1_2/Y DFFSR_208/S
+ AOI21X1
XFILL_17_DFFSR_72 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_28_DFFSR_32 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_0_INVX1_26 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_0_DFFSR_79 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_0_INVX1_164 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_3_AND2X2_31 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_14_DFFSR_120 INVX1_3/gnd DFFSR_23/S FILL
XFILL_7_NAND3X1_97 AND2X2_38/B DFFSR_59/S FILL
XFILL_0_OAI21X1_26 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_28_DFFSR_224 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_18_DFFSR_227 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_4_XOR2X1_9 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_0_NAND3X1_146 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_9_NAND3X1_201 INVX1_1/gnd DFFSR_53/S FILL
XFILL_22_0_0 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_7_OAI22X1_7 AND2X2_38/B DFFSR_59/S FILL
XFILL_5_DFFPOSX1_20 DFFSR_46/gnd DFFSR_62/S FILL
XDFFSR_227 DFFSR_235/D CLKBUF1_21/Y BUFX2_68/Y DFFSR_151/S DFFSR_219/Q BUFX2_7/gnd
+ DFFSR_151/S DFFSR
XFILL_0_DFFSR_117 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_2_NAND2X1_182 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_41_DFFSR_148 INVX1_67/gnd DFFSR_175/S FILL
XFILL_30_4 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_8_DFFSR_86 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_20_2_1 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_25_DFFSR_79 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_36_DFFSR_39 INVX1_3/gnd DFFSR_79/S FILL
XFILL_4_DFFSR_224 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_31_DFFSR_151 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_2_1_0 INVX1_67/gnd DFFSR_201/S FILL
XFILL_45_DFFSR_255 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_21_DFFSR_154 BUFX2_99/A DFFSR_7/S FILL
XFILL_14_DFFPOSX1_39 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_18_4_2 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_35_DFFSR_258 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_3_AOI22X1_10 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_11_DFFSR_157 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_3_NAND2X1_116 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_0_3_1 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_25_DFFSR_261 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_2_AOI22X1_13 AND2X2_38/B DFFSR_23/S FILL
XFILL_6_NOR2X1_33 INVX1_3/gnd DFFSR_23/S FILL
XFILL_15_DFFSR_264 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_1_AOI22X1_16 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_11_OAI22X1_34 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_17_NOR3X1_3 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_10_OAI22X1_37 INVX1_3/gnd DFFSR_23/S FILL
XFILL_0_AOI22X1_19 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_33_DFFSR_86 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_44_DFFSR_46 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_7_DFFSR_151 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_24_DFFPOSX1_28 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_48_DFFSR_182 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_8_NAND3X1_58 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_9_OAI22X1_40 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_38_DFFSR_185 INVX1_39/gnd DFFSR_54/S FILL
XFILL_8_NAND3X1_231 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_17_DFFSR_36 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_0_DFFSR_43 BUFX2_98/A DFFSR_6/S FILL
XFILL_0_INVX1_128 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_7_NAND3X1_61 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_1_DFFSR_261 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_8_OAI22X1_43 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_4_BUFX2_71 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_4_DFFPOSX1_50 INVX1_1/gnd DFFSR_53/S FILL
XFILL_28_DFFSR_188 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_6_NAND3X1_64 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_7_OAI22X1_46 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_18_DFFSR_191 INVX1_67/gnd DFFSR_175/S FILL
XFILL_5_NAND3X1_67 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_6_OAI22X1_49 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_0_NAND3X1_110 XOR2X1_1/gnd DFFSR_151/S FILL
XNAND3X1_64 NOR2X1_27/Y NOR2X1_28/Y NOR2X1_29/Y OR2X2_4/gnd XNOR2X1_4/A DFFSR_32/S
+ NAND3X1
XFILL_10_XOR2X1_6 BUFX2_99/A DFFSR_7/S FILL
XFILL_4_NAND3X1_70 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_5_OAI22X1_52 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_41_DFFSR_93 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_3_NOR2X1_70 XOR2X1_4/gnd DFFSR_91/S FILL
XOAI22X1_49 INVX1_132/Y INVX1_134/Y INVX1_133/Y INVX1_135/Y OR2X2_1/gnd OAI21X1_22/C
+ DFFSR_59/S OAI22X1
XFILL_3_NAND3X1_73 INVX1_1/gnd DFFSR_97/S FILL
XDFFSR_191 DFFSR_183/D CLKBUF1_10/Y BUFX2_64/Y DFFSR_175/S DFFSR_191/D INVX1_67/gnd
+ DFFSR_175/S DFFSR
XFILL_2_NAND2X1_146 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_41_DFFSR_112 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_2_AND2X2_2 BUFX2_99/A DFFSR_7/S FILL
XFILL_2_NAND3X1_76 INVX1_1/gnd DFFSR_53/S FILL
XFILL_8_DFFSR_50 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_25_DFFSR_43 BUFX2_98/A DFFSR_6/S FILL
XFILL_14_DFFSR_83 INVX1_3/gnd DFFSR_79/S FILL
XFILL_4_DFFSR_188 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_31_DFFSR_115 INVX1_1/gnd DFFSR_97/S FILL
XFILL_1_NAND3X1_79 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_45_DFFSR_219 INVX1_67/gnd DFFSR_175/S FILL
XFILL_21_DFFSR_118 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_0_NAND3X1_82 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_35_DFFSR_222 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_0_AND2X2_32 AND2X2_38/B DFFSR_23/S FILL
XFILL_11_DFFSR_121 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_4_NAND2X1_9 BUFX2_79/A DFFSR_6/S FILL
XFILL_25_DFFSR_225 INVX1_67/gnd DFFSR_175/S FILL
XFILL_8_0_2 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_20_DFFSR_5 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_15_DFFSR_228 XOR2X1_1/gnd DFFSR_208/S FILL
XINVX1_84 INVX1_84/A INVX1_39/gnd INVX1_84/Y DFFSR_34/S INVX1
XFILL_44_DFFSR_10 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_33_DFFSR_50 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_5_DFFSR_97 INVX1_1/gnd DFFSR_97/S FILL
XFILL_22_DFFSR_90 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_7_DFFSR_115 INVX1_1/gnd DFFSR_97/S FILL
XFILL_4_OAI22X1_8 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_48_DFFSR_146 BUFX2_79/A DFFSR_7/S FILL
XFILL_4_BUFX2_6 BUFX2_79/A DFFSR_6/S FILL
XFILL_8_NAND3X1_22 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_38_DFFSR_149 BUFX2_72/gnd DFFSR_276/S FILL
XINVX1_202 BUFX2_74/A BUFX2_72/gnd INVX1_202/Y DFFSR_201/S INVX1
XFILL_8_NAND3X1_195 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_1_DFFSR_225 INVX1_67/gnd DFFSR_175/S FILL
XFILL_7_NAND3X1_25 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_4_BUFX2_35 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_28_DFFSR_152 INVX1_1/gnd DFFSR_53/S FILL
XFILL_4_DFFPOSX1_14 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_1_NAND2X1_176 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_6_NAND3X1_28 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_42_DFFSR_256 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_7_OAI22X1_10 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_4_INVX1_199 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_18_DFFSR_155 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_32_DFFSR_259 BUFX2_79/A DFFSR_6/S FILL
XFILL_5_NAND3X1_31 BUFX2_79/A DFFSR_6/S FILL
XFILL_6_OAI22X1_13 INVX1_1/gnd DFFSR_53/S FILL
XFILL_41_DFFSR_1 DFFSR_1/gnd DFFSR_1/S FILL
XNAND3X1_28 NAND3X1_28/A NAND3X1_25/Y AND2X2_9/Y DFFSR_8/gnd NOR2X1_17/A DFFSR_8/S
+ NAND3X1
XFILL_53_4_1 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_22_DFFSR_262 BUFX2_98/A DFFSR_32/S FILL
XFILL_4_NAND3X1_34 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_5_OAI22X1_16 AND2X2_38/B DFFSR_59/S FILL
XFILL_41_DFFSR_57 BUFX2_79/A DFFSR_6/S FILL
XFILL_30_DFFSR_97 INVX1_1/gnd DFFSR_97/S FILL
XFILL_2_INVX1_91 AND2X2_38/B DFFSR_23/S FILL
XFILL_3_NOR2X1_34 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_12_DFFSR_265 INVX1_67/gnd DFFSR_175/S FILL
XOAI22X1_13 INVX1_31/Y OAI22X1_7/B INVX1_32/Y OAI22X1_7/D INVX1_1/gnd NOR2X1_18/B
+ DFFSR_53/S OAI22X1
XFILL_13_DFFPOSX1_33 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_4_OAI22X1_19 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_3_NAND3X1_37 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_2_NAND2X1_110 NOR3X1_6/gnd DFFSR_91/S FILL
XDFFSR_155 INVX1_81/A CLKBUF1_22/Y BUFX2_61/Y DFFSR_59/S DFFSR_155/D OR2X2_1/gnd DFFSR_59/S
+ DFFSR
XFILL_51_6_2 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_2_NAND3X1_40 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_3_OAI22X1_22 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_8_DFFSR_14 INVX1_1/gnd DFFSR_53/S FILL
XFILL_14_DFFSR_47 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_4_DFFSR_152 INVX1_1/gnd DFFSR_53/S FILL
XFILL_1_BUFX2_82 INVX1_1/gnd DFFSR_97/S FILL
XFILL_1_NAND3X1_43 BUFX2_99/A DFFSR_7/S FILL
XFILL_2_OAI22X1_25 INVX1_39/gnd DFFSR_54/S FILL
XFILL_45_DFFSR_183 INVX1_67/gnd DFFSR_175/S FILL
XFILL_0_NAND3X1_46 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_8_DFFSR_259 BUFX2_79/A DFFSR_6/S FILL
XFILL_1_OAI22X1_28 INVX1_3/gnd DFFSR_23/S FILL
XFILL_35_DFFSR_186 BUFX2_99/A DFFSR_92/S FILL
XFILL_23_DFFPOSX1_22 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_0_OAI22X1_31 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_25_DFFSR_189 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_49_DFFSR_64 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_7_NAND3X1_225 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_15_DFFSR_192 INVX1_1/gnd DFFSR_97/S FILL
XFILL_3_DFFPOSX1_44 OR2X2_2/gnd DFFSR_216/S FILL
XINVX1_48 DFFSR_79/Q DFFSR_4/gnd INVX1_48/Y DFFSR_98/S INVX1
XFILL_19_5_0 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_5_DFFSR_61 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_33_DFFSR_14 INVX1_1/gnd DFFSR_53/S FILL
XFILL_11_DFFSR_94 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_22_DFFSR_54 INVX1_39/gnd DFFSR_54/S FILL
XFILL_0_NOR2X1_71 INVX1_1/gnd DFFSR_97/S FILL
XFILL_48_DFFSR_110 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_38_DFFSR_113 BUFX2_99/A DFFSR_92/S FILL
XINVX1_166 AND2X2_36/Y NOR3X1_6/gnd INVX1_166/Y DFFSR_91/S INVX1
XFILL_8_NAND3X1_159 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_1_DFFSR_189 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_28_DFFSR_116 INVX1_3/gnd DFFSR_23/S FILL
XFILL_42_DFFSR_220 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_1_NAND2X1_140 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_7_AND2X2_30 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_18_DFFSR_119 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_32_DFFSR_223 INVX1_39/gnd DFFSR_34/S FILL
XFILL_22_DFFSR_226 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_30_DFFSR_61 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_2_INVX1_55 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_41_DFFSR_21 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_12_DFFSR_229 OR2X2_1/gnd DFFSR_59/S FILL
XDFFSR_119 INVX1_51/A CLKBUF1_5/Y DFFSR_9/R DFFSR_3/S DFFSR_119/D OR2X2_4/gnd DFFSR_3/S
+ DFFSR
XFILL_12_1 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_14_DFFSR_11 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_4_DFFSR_116 INVX1_3/gnd DFFSR_23/S FILL
XFILL_1_BUFX2_46 BUFX2_98/A DFFSR_6/S FILL
XFILL_1_OAI22X1_9 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_45_DFFSR_147 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_0_NAND3X1_10 BUFX2_79/A DFFSR_6/S FILL
XFILL_8_DFFSR_223 INVX1_39/gnd DFFSR_34/S FILL
XFILL_8_DFFSR_4 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_35_DFFSR_150 AND2X2_38/B DFFSR_23/S FILL
XFILL_49_DFFSR_254 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_9_OAI21X1_111 AND2X2_38/B DFFSR_59/S FILL
XFILL_25_DFFSR_153 INVX1_67/gnd DFFSR_201/S FILL
XFILL_1_INVX1_200 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_49_DFFSR_28 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_38_DFFSR_68 BUFX2_98/A DFFSR_6/S FILL
XFILL_39_DFFSR_257 INVX1_39/gnd DFFSR_34/S FILL
XFILL_15_DFFSR_156 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_7_NAND3X1_189 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_29_0_0 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_29_DFFSR_260 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_0_NAND2X1_170 BUFX2_7/gnd DFFSR_216/S FILL
XINVX1_12 DFFSR_82/Q BUFX2_77/gnd INVX1_12/Y DFFSR_5/S INVX1
XDFFSR_65 DFFSR_73/D CLKBUF1_5/Y DFFSR_9/R DFFSR_7/S DFFSR_9/Q BUFX2_79/A DFFSR_7/S
+ DFFSR
XFILL_19_DFFSR_263 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_5_DFFSR_25 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_22_DFFSR_18 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_11_DFFSR_58 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_0_NOR2X1_35 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_27_2_1 INVX1_3/gnd DFFSR_79/S FILL
XFILL_6_OR2X2_4 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_9_1_0 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_8_NAND3X1_123 BUFX2_99/A DFFSR_7/S FILL
XINVX1_130 INVX1_3/A BUFX2_8/gnd INVX1_130/Y DFFSR_51/S INVX1
XFILL_1_DFFSR_153 INVX1_67/gnd DFFSR_201/S FILL
XFILL_4_NOR2X1_6 BUFX2_98/A DFFSR_6/S FILL
XFILL_25_4_2 AND2X2_38/B DFFSR_23/S FILL
XFILL_12_DFFPOSX1_27 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_32_DFFSR_8 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_1_NAND2X1_104 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_42_DFFSR_184 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_4_INVX1_127 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_46_DFFSR_75 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_7_3_1 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_5_DFFSR_260 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_32_DFFSR_187 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_22_DFFSR_190 INVX1_39/gnd DFFSR_34/S FILL
XFILL_2_INVX1_19 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_2_DFFSR_72 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_30_DFFSR_25 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_19_DFFSR_65 BUFX2_79/A DFFSR_7/S FILL
XFILL_5_5_2 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_12_DFFSR_193 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_22_DFFPOSX1_16 INVX1_67/gnd DFFSR_175/S FILL
XFILL_1_BUFX2_10 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_6_NAND3X1_219 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_6_XOR2X1_2 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_45_DFFSR_111 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_2_DFFPOSX1_38 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_8_DFFSR_187 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_35_DFFSR_114 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_49_DFFSR_218 BUFX2_98/A DFFSR_32/S FILL
XAND2X2_34 INVX1_135/A AND2X2_34/B AND2X2_38/B AND2X2_34/Y DFFSR_59/S AND2X2
XFILL_25_DFFSR_117 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_38_DFFSR_32 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_39_DFFSR_221 AND2X2_38/B DFFSR_59/S FILL
XFILL_1_INVX1_164 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_27_DFFSR_72 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_4_AND2X2_31 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_15_DFFSR_120 INVX1_3/gnd DFFSR_23/S FILL
XFILL_7_NAND3X1_153 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_29_DFFSR_224 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_19_DFFSR_227 BUFX2_7/gnd DFFSR_151/S FILL
XDFFSR_29 INVX1_36/A DFFSR_93/CLK DFFSR_5/R DFFSR_5/S DFFSR_5/Q BUFX2_77/gnd DFFSR_5/S
+ DFFSR
XFILL_0_NAND2X1_134 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_11_DFFSR_22 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_8_OAI22X1_7 AND2X2_38/B DFFSR_59/S FILL
XFILL_2_NOR3X1_3 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_1_DFFSR_117 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_17_6 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_34_1 INVX1_1/gnd DFFSR_53/S FILL
XFILL_42_DFFSR_148 INVX1_67/gnd DFFSR_175/S FILL
XFILL_21_DFFPOSX1_46 INVX1_39/gnd DFFSR_34/S FILL
XFILL_35_DFFSR_79 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_46_DFFSR_39 INVX1_3/gnd DFFSR_79/S FILL
XFILL_5_DFFSR_224 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_32_DFFSR_151 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_46_DFFSR_255 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_5_NAND3X1_249 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_22_DFFSR_154 BUFX2_99/A DFFSR_7/S FILL
XFILL_36_DFFSR_258 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_19_DFFSR_29 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_2_DFFSR_36 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_12_DFFSR_157 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_6_BUFX2_64 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_26_DFFSR_261 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_8_OAI21X1_105 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_16_DFFSR_264 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_6_NAND3X1_183 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_20_CLKBUF1_19 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_19_DFFSR_2 BUFX2_79/A DFFSR_7/S FILL
XFILL_43_DFFSR_86 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_19_CLKBUF1_22 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_8_DFFSR_151 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_18_CLKBUF1_25 INVX1_67/gnd DFFSR_201/S FILL
XFILL_49_DFFSR_182 XOR2X1_1/gnd DFFSR_208/S FILL
XNAND3X1_219 AOI21X1_26/Y NAND3X1_219/B NAND3X1_215/Y DFFSR_62/gnd NAND3X1_219/Y DFFSR_62/S
+ NAND3X1
XFILL_17_CLKBUF1_28 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_1_INVX1_128 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_39_DFFSR_185 INVX1_39/gnd DFFSR_54/S FILL
XFILL_27_DFFSR_36 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_16_DFFSR_76 BUFX2_79/A DFFSR_7/S FILL
XFILL_2_DFFSR_261 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_7_NAND3X1_117 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_16_CLKBUF1_31 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_29_DFFSR_188 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_11_DFFPOSX1_21 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_3_BUFX2_3 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_15_CLKBUF1_34 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_19_DFFSR_191 INVX1_67/gnd DFFSR_175/S FILL
XNOR2X1_73 OR2X2_3/B OR2X2_3/A OR2X2_3/gnd NOR2X1_73/Y DFFSR_60/S NOR2X1
XFILL_14_CLKBUF1_37 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_13_CLKBUF1_40 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_4_NOR2X1_70 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_12_CLKBUF1_43 AND2X2_38/B DFFSR_23/S FILL
XFILL_21_DFFPOSX1_10 INVX1_67/gnd DFFSR_201/S FILL
XFILL_42_DFFSR_112 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_11_CLKBUF1_46 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_7_DFFSR_90 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_35_DFFSR_43 BUFX2_98/A DFFSR_6/S FILL
XFILL_24_DFFSR_83 INVX1_3/gnd DFFSR_79/S FILL
XFILL_5_DFFSR_188 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_32_DFFSR_115 INVX1_1/gnd DFFSR_97/S FILL
XFILL_46_DFFSR_219 INVX1_67/gnd DFFSR_175/S FILL
XFILL_10_CLKBUF1_49 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_5_NAND3X1_213 INVX1_39/gnd DFFSR_54/S FILL
XFILL_22_DFFSR_118 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_36_DFFSR_222 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_1_DFFPOSX1_32 INVX1_67/gnd DFFSR_201/S FILL
XFILL_26_5_0 INVX1_3/gnd DFFSR_23/S FILL
XFILL_1_AND2X2_32 AND2X2_38/B DFFSR_23/S FILL
XFILL_12_DFFSR_121 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_6_BUFX2_28 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_5_NAND2X1_9 BUFX2_79/A DFFSR_6/S FILL
XFILL_26_DFFSR_225 INVX1_67/gnd DFFSR_175/S FILL
XFILL_16_DFFSR_228 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_6_NAND3X1_147 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_43_DFFSR_50 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_4_INVX1_84 INVX1_39/gnd DFFSR_34/S FILL
XFILL_6_6_0 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_32_DFFSR_90 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_8_DFFSR_115 INVX1_1/gnd DFFSR_97/S FILL
XFILL_5_OAI22X1_8 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_49_DFFSR_146 BUFX2_79/A DFFSR_7/S FILL
XNAND3X1_183 AOI21X1_28/C AOI21X1_28/B AOI21X1_28/A OR2X2_1/gnd AOI21X1_22/A DFFSR_59/S
+ NAND3X1
XFILL_39_DFFSR_149 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_16_DFFSR_40 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_2_DFFSR_225 INVX1_67/gnd DFFSR_175/S FILL
XFILL_3_BUFX2_75 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_29_DFFSR_152 INVX1_1/gnd DFFSR_53/S FILL
XFILL_43_DFFSR_256 DFFSR_8/gnd DFFSR_60/S FILL
XNAND3X1_2 DFFSR_1/Q NOR2X1_4/Y BUFX2_16/Y BUFX2_99/A AND2X2_6/B DFFSR_7/S NAND3X1
XFILL_20_DFFPOSX1_40 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_19_DFFSR_155 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_33_DFFSR_259 BUFX2_79/A DFFSR_6/S FILL
XNOR2X1_37 NOR2X1_37/A NOR2X1_37/B BUFX2_7/gnd NOR2X1_37/Y DFFSR_216/S NOR2X1
XFILL_23_DFFSR_262 BUFX2_98/A DFFSR_32/S FILL
XFILL_4_NAND3X1_243 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_51_DFFSR_57 BUFX2_79/A DFFSR_6/S FILL
XFILL_40_DFFSR_97 INVX1_1/gnd DFFSR_97/S FILL
XFILL_4_NOR2X1_34 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_13_DFFSR_265 INVX1_67/gnd DFFSR_175/S FILL
XFILL_1_AND2X2_6 BUFX2_99/A DFFSR_7/S FILL
XFILL_11_CLKBUF1_10 INVX1_67/gnd DFFSR_201/S FILL
XFILL_24_DFFSR_47 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_7_DFFSR_54 INVX1_39/gnd DFFSR_54/S FILL
XFILL_13_DFFSR_87 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_5_DFFSR_152 INVX1_1/gnd DFFSR_53/S FILL
XFILL_46_DFFSR_183 INVX1_67/gnd DFFSR_175/S FILL
XFILL_10_CLKBUF1_13 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_36_0_0 BUFX2_99/A DFFSR_92/S FILL
XFILL_5_NAND3X1_177 AND2X2_38/B DFFSR_59/S FILL
XFILL_9_DFFSR_259 BUFX2_79/A DFFSR_6/S FILL
XFILL_36_DFFSR_186 BUFX2_99/A DFFSR_92/S FILL
XFILL_9_CLKBUF1_16 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_34_2_1 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_26_DFFSR_189 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_7_DFFSR_1 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_10_DFFSR_9 BUFX2_79/A DFFSR_6/S FILL
XFILL_16_DFFSR_192 INVX1_1/gnd DFFSR_97/S FILL
XFILL_8_CLKBUF1_19 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_6_NAND3X1_111 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_32_4_2 INVX1_1/gnd DFFSR_97/S FILL
XFILL_7_CLKBUF1_22 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_10_DFFPOSX1_15 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_4_INVX1_48 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_43_DFFSR_14 INVX1_1/gnd DFFSR_53/S FILL
XFILL_21_DFFSR_94 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_32_DFFSR_54 INVX1_39/gnd DFFSR_54/S FILL
XFILL_6_CLKBUF1_25 INVX1_67/gnd DFFSR_201/S FILL
XFILL_1_NOR2X1_71 INVX1_1/gnd DFFSR_97/S FILL
XFILL_49_DFFSR_110 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_5_CLKBUF1_28 OR2X2_4/gnd DFFSR_3/S FILL
XNAND3X1_147 INVX1_144/Y OAI21X1_32/Y OAI21X1_33/Y OR2X2_1/gnd AOI21X1_14/B DFFSR_51/S
+ NAND3X1
XFILL_39_DFFSR_113 BUFX2_99/A DFFSR_92/S FILL
XCLKBUF1_25 BUFX2_3/Y INVX1_67/gnd CLKBUF1_25/Y DFFSR_201/S CLKBUF1
XFILL_4_CLKBUF1_31 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_5_OR2X2_1 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_2_DFFSR_189 BUFX2_8/gnd DFFSR_51/S FILL
XOR2X2_5 OR2X2_5/A OR2X2_5/B BUFX2_8/gnd OR2X2_5/Y DFFSR_81/S OR2X2
XFILL_3_BUFX2_39 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_29_DFFSR_116 INVX1_3/gnd DFFSR_23/S FILL
XFILL_3_CLKBUF1_34 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_43_DFFSR_220 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_8_AND2X2_30 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_19_DFFSR_119 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_2_CLKBUF1_37 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_33_DFFSR_223 INVX1_39/gnd DFFSR_34/S FILL
XFILL_31_DFFSR_5 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_23_DFFSR_226 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_4_NAND3X1_207 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_1_CLKBUF1_40 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_1_INVX1_95 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_40_DFFSR_61 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_51_DFFSR_21 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_13_DFFSR_229 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_0_DFFPOSX1_26 AND2X2_38/B DFFSR_23/S FILL
XFILL_0_CLKBUF1_43 AND2X2_38/B DFFSR_23/S FILL
XFILL_7_DFFSR_18 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_24_DFFSR_11 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_5_DFFSR_116 INVX1_3/gnd DFFSR_23/S FILL
XFILL_13_DFFSR_51 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_0_BUFX2_86 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_2_OAI22X1_9 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_46_DFFSR_147 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_5_NAND3X1_141 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_9_DFFSR_223 INVX1_39/gnd DFFSR_34/S FILL
XFILL_36_DFFSR_150 AND2X2_38/B DFFSR_23/S FILL
XFILL_50_DFFSR_254 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_26_DFFSR_153 INVX1_67/gnd DFFSR_201/S FILL
XFILL_2_INVX1_200 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_40_DFFSR_257 INVX1_39/gnd DFFSR_34/S FILL
XFILL_48_DFFSR_68 BUFX2_98/A DFFSR_6/S FILL
XFILL_16_DFFSR_156 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_30_DFFSR_260 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_20_DFFSR_263 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_4_DFFSR_65 BUFX2_79/A DFFSR_7/S FILL
XFILL_19_DFFPOSX1_34 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_21_DFFSR_58 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_10_DFFSR_98 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_32_DFFSR_18 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_1_NOR2X1_35 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_10_DFFSR_266 INVX1_67/gnd DFFSR_201/S FILL
XNAND3X1_111 NAND3X1_111/A NAND3X1_110/Y AOI22X1_14/Y XOR2X1_1/gnd NOR2X1_52/B DFFSR_151/S
+ NAND3X1
XFILL_3_NAND3X1_237 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_2_DFFSR_153 INVX1_67/gnd DFFSR_201/S FILL
XFILL_43_DFFSR_184 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_6_DFFSR_260 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_33_DFFSR_187 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_4_NAND3X1_171 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_23_DFFSR_190 INVX1_39/gnd DFFSR_34/S FILL
XFILL_40_DFFSR_25 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_29_DFFSR_65 BUFX2_79/A DFFSR_7/S FILL
XFILL_1_INVX1_59 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_13_DFFSR_193 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_9_DFFPOSX1_45 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_13_DFFSR_15 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_0_BUFX2_50 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_46_DFFSR_111 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_5_NAND3X1_105 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_9_DFFSR_187 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_36_DFFSR_114 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_50_DFFSR_218 BUFX2_98/A DFFSR_32/S FILL
XFILL_26_DFFSR_117 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_48_DFFSR_32 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_40_DFFSR_221 AND2X2_38/B DFFSR_59/S FILL
XFILL_2_INVX1_164 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_37_DFFSR_72 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_5_AND2X2_31 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_16_DFFSR_120 INVX1_3/gnd DFFSR_23/S FILL
XFILL_30_DFFSR_224 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_20_DFFSR_227 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_4_DFFSR_29 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_21_DFFSR_22 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_10_DFFSR_62 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_10_DFFSR_230 INVX1_67/gnd DFFSR_201/S FILL
XFILL_3_NAND3X1_201 INVX1_1/gnd DFFSR_53/S FILL
XFILL_9_OAI22X1_7 AND2X2_38/B DFFSR_59/S FILL
XFILL_2_DFFSR_117 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_33_5_0 INVX1_1/gnd DFFSR_53/S FILL
XFILL_43_DFFSR_148 INVX1_67/gnd DFFSR_175/S FILL
XFILL_45_DFFSR_79 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_6_DFFSR_224 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_33_DFFSR_151 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_47_DFFSR_255 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_23_DFFSR_154 BUFX2_99/A DFFSR_7/S FILL
XFILL_4_NAND3X1_135 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_37_DFFSR_258 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_29_DFFSR_29 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_1_DFFSR_76 BUFX2_79/A DFFSR_7/S FILL
XFILL_1_INVX1_23 BUFX2_99/A DFFSR_7/S FILL
XFILL_18_DFFSR_69 BUFX2_98/A DFFSR_32/S FILL
XFILL_13_DFFSR_157 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_27_DFFSR_261 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_6_NAND2X1_171 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_17_DFFSR_264 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_22_DFFPOSX1_1 INVX1_39/gnd DFFSR_34/S FILL
XFILL_0_BUFX2_14 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_5_XOR2X1_6 BUFX2_99/A DFFSR_7/S FILL
XFILL_21_DFFPOSX1_4 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_9_DFFSR_151 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_43_DFFSR_8 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_20_DFFPOSX1_7 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_18_DFFPOSX1_28 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_50_DFFSR_182 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_9_DFFSR_83 INVX1_3/gnd DFFSR_79/S FILL
XFILL_2_INVX1_128 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_40_DFFSR_185 INVX1_39/gnd DFFSR_54/S FILL
XFILL_37_DFFSR_36 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_26_DFFSR_76 BUFX2_79/A DFFSR_7/S FILL
XFILL_2_NAND3X1_231 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_3_DFFSR_261 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_30_DFFSR_188 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_20_DFFSR_191 INVX1_67/gnd DFFSR_175/S FILL
XFILL_10_DFFSR_26 BUFX2_79/A DFFSR_6/S FILL
XFILL_10_DFFSR_194 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_43_0_0 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_5_NOR2X1_70 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_3_NAND3X1_165 INVX1_39/gnd DFFSR_34/S FILL
XFILL_43_DFFSR_112 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_8_DFFPOSX1_39 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_41_2_1 BUFX2_98/A DFFSR_32/S FILL
XFILL_45_DFFSR_43 BUFX2_98/A DFFSR_6/S FILL
XFILL_34_DFFSR_83 INVX1_3/gnd DFFSR_79/S FILL
XFILL_6_DFFSR_188 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_33_DFFSR_115 INVX1_1/gnd DFFSR_97/S FILL
XFILL_47_DFFSR_219 INVX1_67/gnd DFFSR_175/S FILL
XFILL_23_DFFSR_118 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_37_DFFSR_222 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_1_DFFSR_40 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_39_4_2 BUFX2_79/A DFFSR_6/S FILL
XFILL_18_DFFSR_33 BUFX2_98/A DFFSR_32/S FILL
XFILL_2_AND2X2_32 AND2X2_38/B DFFSR_23/S FILL
XFILL_13_DFFSR_121 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_6_NAND2X1_9 BUFX2_79/A DFFSR_6/S FILL
XFILL_5_BUFX2_68 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_27_DFFSR_225 INVX1_67/gnd DFFSR_175/S FILL
XFILL_6_NAND2X1_135 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_17_DFFSR_228 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_11_XOR2X1_3 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_42_DFFSR_90 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_9_DFFSR_115 INVX1_1/gnd DFFSR_97/S FILL
XNAND2X1_171 INVX1_209/Y NOR3X1_6/C NOR3X1_6/gnd NOR2X1_76/B DFFSR_79/S NAND2X1
XFILL_6_OAI22X1_8 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_50_DFFSR_146 BUFX2_79/A DFFSR_7/S FILL
XFILL_4_OAI21X1_117 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_27_DFFPOSX1_47 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_8_AOI21X1_63 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_40_DFFSR_149 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_9_DFFSR_47 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_26_DFFSR_40 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_15_DFFSR_80 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_7_AOI21X1_66 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_3_DFFSR_225 INVX1_67/gnd DFFSR_175/S FILL
XFILL_2_NAND3X1_195 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_30_DFFSR_152 INVX1_1/gnd DFFSR_53/S FILL
XFILL_6_AOI21X1_69 INVX1_1/gnd DFFSR_97/S FILL
XFILL_44_DFFSR_256 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_20_DFFSR_155 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_34_DFFSR_259 BUFX2_79/A DFFSR_6/S FILL
XAOI21X1_69 XOR2X1_14/Y NOR2X1_81/Y BUFX2_40/Y INVX1_1/gnd AOI21X1_69/Y DFFSR_97/S
+ AOI21X1
XFILL_10_DFFSR_158 INVX1_3/gnd DFFSR_23/S FILL
XFILL_24_DFFSR_262 BUFX2_98/A DFFSR_32/S FILL
XFILL_50_DFFSR_97 INVX1_1/gnd DFFSR_97/S FILL
XFILL_5_NOR2X1_34 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_3_NAND3X1_129 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_30_DFFSR_2 BUFX2_79/A DFFSR_7/S FILL
XFILL_14_DFFSR_265 INVX1_67/gnd DFFSR_175/S FILL
XFILL_34_DFFSR_47 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_6_DFFSR_94 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_5_NAND2X1_165 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_23_DFFSR_87 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_6_DFFSR_152 INVX1_1/gnd DFFSR_53/S FILL
XFILL_47_DFFSR_183 INVX1_67/gnd DFFSR_175/S FILL
XFILL_37_DFFSR_186 BUFX2_99/A DFFSR_92/S FILL
XBUFX2_72 BUFX2_72/A BUFX2_72/gnd dout[1] DFFSR_201/S BUFX2
XFILL_0_DFFSR_262 BUFX2_98/A DFFSR_32/S FILL
XFILL_5_BUFX2_32 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_10_DFFPOSX1_1 INVX1_39/gnd DFFSR_34/S FILL
XFILL_27_DFFSR_189 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_17_DFFPOSX1_22 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_17_DFFSR_192 INVX1_1/gnd DFFSR_97/S FILL
XFILL_1_NAND3X1_225 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_9_DFFPOSX1_4 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_3_INVX1_88 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_8_DFFPOSX1_7 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_31_DFFSR_94 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_42_DFFSR_54 INVX1_39/gnd DFFSR_54/S FILL
XFILL_9_AOI21X1_24 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_2_NOR2X1_71 INVX1_1/gnd DFFSR_97/S FILL
XNAND2X1_135 DFFSR_34/S INVX1_193/A DFFSR_34/gnd OAI21X1_104/C DFFSR_34/S NAND2X1
XFILL_50_DFFSR_110 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_8_AOI21X1_27 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_27_DFFPOSX1_11 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_40_DFFSR_113 BUFX2_99/A DFFSR_92/S FILL
XFILL_9_DFFSR_11 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_15_DFFSR_44 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_7_AOI21X1_30 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_2_NAND3X1_159 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_3_DFFSR_189 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_2_BUFX2_79 BUFX2_79/A DFFSR_7/S FILL
XFILL_30_DFFSR_116 INVX1_3/gnd DFFSR_23/S FILL
XFILL_15_0_1 INVX1_39/gnd DFFSR_34/S FILL
XFILL_6_AOI21X1_33 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_44_DFFSR_220 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_20_DFFSR_119 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_7_DFFPOSX1_33 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_5_AOI21X1_36 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_34_DFFSR_223 INVX1_39/gnd DFFSR_34/S FILL
XFILL_10_DFFSR_122 BUFX2_79/A DFFSR_7/S FILL
XAOI21X1_33 INVX1_157/Y OAI21X1_52/Y AOI21X1_33/C XOR2X1_1/gnd AOI21X1_33/Y DFFSR_208/S
+ AOI21X1
XFILL_13_2_2 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_4_AOI21X1_39 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_24_DFFSR_226 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_50_DFFSR_61 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_0_AOI21X1_1 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_3_AOI21X1_42 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_14_DFFSR_229 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_2_AOI21X1_45 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_6_DFFSR_58 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_34_DFFSR_11 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_5_NAND2X1_129 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_12_DFFSR_91 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_6_DFFSR_116 INVX1_3/gnd DFFSR_23/S FILL
XFILL_23_DFFSR_51 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_1_AOI21X1_48 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_3_OAI22X1_9 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_47_DFFSR_147 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_0_AOI21X1_51 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_37_DFFSR_150 AND2X2_38/B DFFSR_23/S FILL
XBUFX2_36 rst OR2X2_2/gnd BUFX2_36/Y DFFSR_175/S BUFX2
XFILL_51_DFFSR_254 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_0_DFFSR_226 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_27_DFFSR_153 INVX1_67/gnd DFFSR_201/S FILL
XFILL_3_OAI21X1_111 AND2X2_38/B DFFSR_59/S FILL
XFILL_3_INVX1_200 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_26_DFFPOSX1_41 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_41_DFFSR_257 INVX1_39/gnd DFFSR_34/S FILL
XFILL_17_DFFSR_156 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_31_DFFSR_260 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_8_OAI21X1_75 INVX1_39/gnd DFFSR_54/S FILL
XFILL_1_NAND3X1_189 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_7_OAI21X1_78 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_6_NAND2X1_96 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_40_5_0 BUFX2_98/A DFFSR_6/S FILL
XFILL_21_DFFSR_263 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_31_DFFSR_58 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_3_INVX1_52 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_20_DFFSR_98 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_42_DFFSR_18 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_2_NOR2X1_35 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_6_OAI21X1_81 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_5_NAND2X1_99 INVX1_39/gnd DFFSR_54/S FILL
XFILL_11_DFFSR_266 INVX1_67/gnd DFFSR_201/S FILL
XNAND2X1_96 INVX1_175/A AND2X2_33/B OR2X2_6/gnd INVX1_167/A DFFSR_53/S NAND2X1
XFILL_5_OAI21X1_84 BUFX2_98/A DFFSR_6/S FILL
XOAI21X1_81 OAI21X1_80/A OAI21X1_80/B INVX1_179/Y OR2X2_3/gnd AOI21X1_39/A DFFSR_4/S
+ OAI21X1
XFILL_3_DFFSR_153 INVX1_67/gnd DFFSR_201/S FILL
XFILL_2_NAND3X1_123 BUFX2_99/A DFFSR_7/S FILL
XFILL_4_OAI21X1_87 BUFX2_79/A DFFSR_7/S FILL
XFILL_2_BUFX2_43 AND2X2_38/B DFFSR_23/S FILL
XFILL_44_DFFSR_184 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_3_OAI21X1_90 BUFX2_98/A DFFSR_32/S FILL
XFILL_7_DFFSR_260 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_4_NAND2X1_159 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_34_DFFSR_187 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_2_OAI21X1_93 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_21_DFFSR_9 BUFX2_79/A DFFSR_6/S FILL
XFILL_24_DFFSR_190 INVX1_39/gnd DFFSR_34/S FILL
XFILL_50_DFFSR_25 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_1_OAI21X1_96 AND2X2_38/B DFFSR_59/S FILL
XFILL_0_INVX1_99 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_39_DFFSR_65 BUFX2_79/A DFFSR_7/S FILL
XFILL_14_DFFSR_193 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_0_OAI21X1_99 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_16_DFFPOSX1_16 INVX1_67/gnd DFFSR_175/S FILL
XFILL_6_DFFSR_22 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_23_DFFSR_15 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_12_DFFSR_55 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_1_AOI21X1_12 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_47_DFFSR_111 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_0_NAND3X1_219 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_0_AOI21X1_15 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_37_DFFSR_114 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_5_NOR2X1_3 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_0_DFFSR_190 INVX1_39/gnd DFFSR_34/S FILL
XFILL_27_DFFSR_117 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_42_DFFSR_5 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_41_DFFSR_221 AND2X2_38/B DFFSR_59/S FILL
XFILL_3_INVX1_164 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_47_DFFSR_72 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_6_AND2X2_31 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_17_DFFSR_120 INVX1_3/gnd DFFSR_23/S FILL
XFILL_50_0_0 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_31_DFFSR_224 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_8_OAI21X1_39 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_1_NAND3X1_153 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_21_DFFSR_227 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_7_OAI21X1_42 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_6_NAND2X1_60 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_31_DFFSR_22 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_3_DFFSR_69 BUFX2_98/A DFFSR_32/S FILL
XFILL_3_INVX1_16 BUFX2_99/A DFFSR_7/S FILL
XFILL_20_DFFSR_62 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_6_DFFPOSX1_27 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_48_2_1 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_5_NAND2X1_63 AND2X2_38/B DFFSR_59/S FILL
XFILL_6_OAI21X1_45 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_11_DFFSR_230 INVX1_67/gnd DFFSR_201/S FILL
XNAND2X1_60 AND2X2_35/A INVX1_135/A DFFSR_34/gnd NOR2X1_66/B DFFSR_34/S NAND2X1
XFILL_5_OAI21X1_48 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_4_NAND2X1_66 BUFX2_8/gnd DFFSR_81/S FILL
XOAI21X1_45 INVX1_131/Y NAND2X1_79/Y OAI21X1_45/C DFFSR_62/gnd OAI21X1_45/Y DFFSR_208/S
+ OAI21X1
XFILL_3_DFFSR_117 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_46_4_2 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_3_NAND2X1_69 INVX1_3/gnd DFFSR_23/S FILL
XFILL_4_OAI21X1_51 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_44_DFFSR_148 INVX1_67/gnd DFFSR_175/S FILL
XFILL_2_NAND2X1_72 AND2X2_38/B DFFSR_59/S FILL
XFILL_15_DFFPOSX1_46 INVX1_39/gnd DFFSR_34/S FILL
XFILL_3_OAI21X1_54 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_7_DFFSR_224 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_34_DFFSR_151 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_4_NAND2X1_123 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_1_NAND2X1_75 INVX1_3/gnd DFFSR_79/S FILL
XFILL_2_OAI21X1_57 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_48_DFFSR_255 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_11_AOI22X1_23 INVX1_39/gnd DFFSR_34/S FILL
XFILL_24_DFFSR_154 BUFX2_99/A DFFSR_7/S FILL
XFILL_0_NAND2X1_78 AND2X2_38/B DFFSR_23/S FILL
XFILL_38_DFFSR_258 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_39_DFFSR_29 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_0_INVX1_201 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_0_INVX1_63 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_1_OAI21X1_60 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_28_DFFSR_69 BUFX2_98/A DFFSR_32/S FILL
XFILL_10_AOI22X1_26 INVX1_1/gnd DFFSR_97/S FILL
XFILL_14_DFFSR_157 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_28_DFFSR_261 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_0_OAI21X1_63 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_2_OAI21X1_105 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_18_DFFSR_264 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_9_AOI22X1_29 INVX1_1/gnd DFFSR_53/S FILL
XFILL_25_DFFPOSX1_35 INVX1_39/gnd DFFSR_54/S FILL
XFILL_12_DFFSR_19 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_0_NAND3X1_183 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_14_3_0 INVX1_39/gnd DFFSR_54/S FILL
XNOR2X1_7 OR2X2_1/A BUFX2_7/Y BUFX2_98/A NOR2X1_7/Y DFFSR_32/S NOR2X1
XFILL_51_DFFSR_182 XOR2X1_1/gnd DFFSR_208/S FILL
XDFFSR_264 DFFSR_8/D CLKBUF1_4/Y DFFSR_257/R DFFSR_264/S DFFSR_264/D DFFSR_4/gnd DFFSR_98/S
+ DFFSR
XFILL_0_DFFSR_154 BUFX2_99/A DFFSR_7/S FILL
XFILL_12_5_1 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_3_INVX1_128 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_41_DFFSR_185 INVX1_39/gnd DFFSR_54/S FILL
XFILL_47_DFFSR_36 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_36_DFFSR_76 BUFX2_79/A DFFSR_7/S FILL
XFILL_4_DFFSR_261 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_31_DFFSR_188 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_1_NAND3X1_117 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_21_DFFSR_191 INVX1_67/gnd DFFSR_175/S FILL
XFILL_6_NAND2X1_24 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_3_DFFSR_33 BUFX2_98/A DFFSR_32/S FILL
XFILL_20_DFFSR_26 BUFX2_79/A DFFSR_6/S FILL
XFILL_3_NAND2X1_153 BUFX2_98/A DFFSR_32/S FILL
XFILL_5_NAND2X1_27 AND2X2_38/B DFFSR_23/S FILL
XFILL_11_DFFSR_194 DFFSR_1/gnd DFFSR_81/S FILL
XNAND2X1_24 DFFSR_39/Q AND2X2_5/Y OR2X2_3/gnd NAND3X1_52/A DFFSR_4/S NAND2X1
XFILL_4_NAND2X1_30 AND2X2_38/B DFFSR_23/S FILL
XFILL_5_OAI21X1_12 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_6_NOR2X1_70 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_8_4 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_9_DFFSR_8 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_3_NAND2X1_33 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_4_OAI21X1_15 INVX1_3/gnd DFFSR_79/S FILL
XDFFPOSX1_27 NAND2X1_149/B CLKBUF1_49/Y AOI21X1_51/Y DFFSR_34/gnd DFFSR_1/S DFFPOSX1
XFILL_44_DFFSR_112 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_15_DFFPOSX1_10 INVX1_67/gnd DFFSR_201/S FILL
XFILL_2_NAND2X1_36 INVX1_3/gnd DFFSR_79/S FILL
XFILL_3_OAI21X1_18 INVX1_39/gnd DFFSR_34/S FILL
XFILL_44_DFFSR_83 INVX1_3/gnd DFFSR_79/S FILL
XFILL_7_DFFSR_188 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_34_DFFSR_115 INVX1_1/gnd DFFSR_97/S FILL
XFILL_1_NAND2X1_39 BUFX2_98/A DFFSR_6/S FILL
XFILL_2_OAI21X1_21 AND2X2_38/B DFFSR_59/S FILL
XFILL_48_DFFSR_219 INVX1_67/gnd DFFSR_175/S FILL
XFILL_24_DFFSR_118 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_0_NAND2X1_42 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_8_NAND3X1_95 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_38_DFFSR_222 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_0_INVX1_27 BUFX2_99/A DFFSR_7/S FILL
XFILL_0_INVX1_165 BUFX2_99/A DFFSR_92/S FILL
XFILL_1_OAI21X1_24 DFFSR_34/gnd DFFSR_1/S FILL
XAOI21X1_3 AND2X2_27/B AOI21X1_3/B BUFX2_38/Y DFFSR_34/gnd AOI21X1_3/Y DFFSR_1/S AOI21X1
XFILL_0_DFFSR_80 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_28_DFFSR_33 BUFX2_98/A DFFSR_32/S FILL
XFILL_3_AND2X2_32 AND2X2_38/B DFFSR_23/S FILL
XFILL_17_DFFSR_73 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_14_DFFSR_121 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_7_NAND3X1_98 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_28_DFFSR_225 INVX1_67/gnd DFFSR_175/S FILL
XFILL_0_OAI21X1_27 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_18_DFFSR_228 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_0_NAND3X1_147 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_22_0_1 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_9_NAND3X1_202 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_7_OAI22X1_8 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_5_DFFPOSX1_21 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_0_DFFSR_118 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_51_DFFSR_146 BUFX2_79/A DFFSR_7/S FILL
XDFFSR_228 DFFSR_228/Q CLKBUF1_21/Y BUFX2_68/Y DFFSR_208/S DFFSR_220/Q XOR2X1_1/gnd
+ DFFSR_208/S DFFSR
XFILL_41_DFFSR_149 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_30_5 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_36_DFFSR_40 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_8_DFFSR_87 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_20_2_2 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_25_DFFSR_80 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_4_DFFSR_225 INVX1_67/gnd DFFSR_175/S FILL
XFILL_31_DFFSR_152 INVX1_1/gnd DFFSR_53/S FILL
XFILL_2_1_1 INVX1_67/gnd DFFSR_201/S FILL
XFILL_45_DFFSR_256 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_21_DFFSR_155 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_35_DFFSR_259 BUFX2_79/A DFFSR_6/S FILL
XFILL_14_DFFPOSX1_40 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_3_AOI22X1_11 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_3_NAND2X1_117 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_11_DFFSR_158 INVX1_3/gnd DFFSR_23/S FILL
XFILL_0_3_2 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_2_AOI22X1_14 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_25_DFFSR_262 BUFX2_98/A DFFSR_32/S FILL
XINVX1_1 INVX1_1/A INVX1_1/gnd INVX1_1/Y DFFSR_53/S INVX1
XFILL_6_NOR2X1_34 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_15_DFFSR_265 INVX1_67/gnd DFFSR_175/S FILL
XFILL_11_OAI22X1_35 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_17_NOR3X1_4 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_1_AOI22X1_17 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_10_OAI22X1_38 AND2X2_38/B DFFSR_23/S FILL
XFILL_0_AOI22X1_20 INVX1_39/gnd DFFSR_34/S FILL
XFILL_33_DFFSR_87 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_44_DFFSR_47 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_7_DFFSR_152 INVX1_1/gnd DFFSR_53/S FILL
XFILL_24_DFFPOSX1_29 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_48_DFFSR_183 INVX1_67/gnd DFFSR_175/S FILL
XFILL_8_NAND3X1_59 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_9_OAI22X1_41 INVX1_39/gnd DFFSR_54/S FILL
XFILL_0_DFFSR_44 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_8_NAND3X1_232 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_38_DFFSR_186 BUFX2_99/A DFFSR_92/S FILL
XFILL_0_INVX1_129 AND2X2_38/B DFFSR_23/S FILL
XFILL_17_DFFSR_37 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_4_BUFX2_72 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_47_5_0 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_7_NAND3X1_62 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_1_DFFSR_262 BUFX2_98/A DFFSR_32/S FILL
XFILL_8_OAI22X1_44 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_28_DFFSR_189 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_7_OAI22X1_47 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_6_NAND3X1_65 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_18_DFFSR_192 INVX1_1/gnd DFFSR_97/S FILL
XFILL_5_NAND3X1_68 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_6_OAI22X1_50 INVX1_3/gnd DFFSR_23/S FILL
XFILL_0_NAND3X1_111 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_10_XOR2X1_7 BUFX2_98/A DFFSR_6/S FILL
XNAND3X1_65 DFFSR_169/Q BUFX2_27/Y BUFX2_23/Y DFFSR_62/gnd NAND3X1_68/B DFFSR_208/S
+ NAND3X1
XFILL_4_NAND3X1_71 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_41_DFFSR_94 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_3_NOR2X1_71 INVX1_1/gnd DFFSR_97/S FILL
XOAI22X1_50 OAI21X1_31/C NOR2X1_70/A INVX1_151/A OAI22X1_50/D INVX1_3/gnd AOI21X1_28/C
+ DFFSR_23/S OAI22X1
XFILL_3_NAND3X1_74 INVX1_1/gnd DFFSR_97/S FILL
XFILL_2_NAND2X1_147 OR2X2_2/gnd DFFSR_216/S FILL
XDFFSR_192 DFFSR_184/D CLKBUF1_39/Y BUFX2_63/Y DFFSR_97/S DFFSR_192/D INVX1_1/gnd
+ DFFSR_97/S DFFSR
XFILL_2_AND2X2_3 INVX1_1/gnd DFFSR_53/S FILL
XFILL_2_NAND3X1_77 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_41_DFFSR_113 BUFX2_99/A DFFSR_92/S FILL
XFILL_25_DFFSR_44 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_8_DFFSR_51 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_14_DFFSR_84 BUFX2_99/A DFFSR_7/S FILL
XFILL_4_DFFSR_189 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_1_NAND3X1_80 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_31_DFFSR_116 INVX1_3/gnd DFFSR_23/S FILL
XFILL_45_DFFSR_220 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_21_DFFSR_119 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_0_NAND3X1_83 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_35_DFFSR_223 INVX1_39/gnd DFFSR_34/S FILL
XFILL_0_AND2X2_33 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_11_DFFSR_122 BUFX2_79/A DFFSR_7/S FILL
XFILL_25_DFFSR_226 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_1_AOI21X1_1 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_20_DFFSR_6 BUFX2_79/A DFFSR_6/S FILL
XFILL_15_DFFSR_229 OR2X2_1/gnd DFFSR_59/S FILL
XINVX1_85 INVX1_85/A DFFSR_46/gnd INVX1_85/Y DFFSR_54/S INVX1
XFILL_5_DFFSR_98 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_22_DFFSR_91 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_7_DFFSR_116 INVX1_3/gnd DFFSR_23/S FILL
XFILL_33_DFFSR_51 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_44_DFFSR_11 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_9_NAND3X1_20 BUFX2_99/A DFFSR_7/S FILL
XFILL_4_OAI22X1_9 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_48_DFFSR_147 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_8_NAND3X1_23 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_4_BUFX2_7 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_38_DFFSR_150 AND2X2_38/B DFFSR_23/S FILL
XFILL_8_NAND3X1_196 DFFSR_46/gnd DFFSR_62/S FILL
XINVX1_203 BUFX2_75/A BUFX2_72/gnd INVX1_203/Y DFFSR_276/S INVX1
XFILL_4_BUFX2_36 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_7_NAND3X1_26 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_1_DFFSR_226 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_4_DFFPOSX1_15 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_28_DFFSR_153 INVX1_67/gnd DFFSR_201/S FILL
XFILL_1_NAND2X1_177 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_42_DFFSR_257 INVX1_39/gnd DFFSR_34/S FILL
XFILL_4_INVX1_200 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_6_NAND3X1_29 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_7_OAI22X1_11 BUFX2_99/A DFFSR_92/S FILL
XFILL_18_DFFSR_156 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_32_DFFSR_260 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_6_OAI22X1_14 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_5_NAND3X1_32 BUFX2_79/A DFFSR_7/S FILL
XFILL_41_DFFSR_2 BUFX2_79/A DFFSR_7/S FILL
XNAND3X1_29 DFFSR_68/D BUFX2_21/Y BUFX2_12/Y OR2X2_4/gnd NAND3X1_31/A DFFSR_32/S NAND3X1
XFILL_4_NAND3X1_35 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_53_4_2 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_22_DFFSR_263 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_9_NAND3X1_130 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_41_DFFSR_58 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_5_OAI22X1_17 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_2_INVX1_92 AND2X2_38/B DFFSR_23/S FILL
XFILL_3_NOR2X1_35 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_30_DFFSR_98 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_13_DFFPOSX1_34 OR2X2_2/gnd DFFSR_216/S FILL
XOAI22X1_14 INVX1_33/Y OAI22X1_2/B INVX1_34/Y OAI22X1_2/D OR2X2_4/gnd NOR2X1_18/A
+ DFFSR_3/S OAI22X1
XFILL_12_DFFSR_266 INVX1_67/gnd DFFSR_201/S FILL
XFILL_4_OAI22X1_20 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_3_NAND3X1_38 BUFX2_98/A DFFSR_32/S FILL
XDFFSR_156 INVX1_88/A CLKBUF1_2/Y BUFX2_67/Y DFFSR_175/S DFFSR_156/D OR2X2_2/gnd DFFSR_175/S
+ DFFSR
XFILL_2_NAND2X1_111 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_3_OAI22X1_23 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_2_NAND3X1_41 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_8_DFFSR_15 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_14_DFFSR_48 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_4_DFFSR_153 INVX1_67/gnd DFFSR_201/S FILL
XFILL_1_BUFX2_83 BUFX2_79/A DFFSR_7/S FILL
XFILL_1_NAND3X1_44 BUFX2_99/A DFFSR_7/S FILL
XFILL_2_OAI22X1_26 INVX1_39/gnd DFFSR_54/S FILL
XFILL_45_DFFSR_184 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_0_NAND3X1_47 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_8_DFFSR_260 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_1_OAI22X1_29 INVX1_3/gnd DFFSR_79/S FILL
XFILL_35_DFFSR_187 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_23_DFFPOSX1_23 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_0_OAI22X1_32 INVX1_39/gnd DFFSR_54/S FILL
XFILL_25_DFFSR_190 INVX1_39/gnd DFFSR_34/S FILL
XFILL_21_3_0 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_49_DFFSR_65 BUFX2_79/A DFFSR_7/S FILL
XFILL_15_DFFSR_193 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_7_NAND3X1_226 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_3_DFFPOSX1_45 OR2X2_1/gnd DFFSR_59/S FILL
XINVX1_49 DFFSR_23/Q OR2X2_6/gnd INVX1_49/Y DFFSR_53/S INVX1
XFILL_19_5_1 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_33_DFFSR_15 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_22_DFFSR_55 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_11_DFFSR_95 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_5_DFFSR_62 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_0_NOR2X1_72 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_1_4_0 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_48_DFFSR_111 DFFSR_8/gnd DFFSR_8/S FILL
XINVX1_167 INVX1_167/A OR2X2_6/gnd INVX1_167/Y DFFSR_53/S INVX1
XFILL_38_DFFSR_114 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_8_NAND3X1_160 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_1_DFFSR_190 INVX1_39/gnd DFFSR_34/S FILL
XFILL_28_DFFSR_117 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_42_DFFSR_221 AND2X2_38/B DFFSR_59/S FILL
XFILL_4_INVX1_164 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_1_NAND2X1_141 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_7_AND2X2_31 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_18_DFFSR_120 INVX1_3/gnd DFFSR_23/S FILL
XFILL_32_DFFSR_224 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_22_DFFSR_227 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_41_DFFSR_22 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_2_INVX1_56 BUFX2_98/A DFFSR_6/S FILL
XFILL_30_DFFSR_62 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_12_DFFSR_230 INVX1_67/gnd DFFSR_201/S FILL
XDFFSR_120 INVX1_58/A CLKBUF1_18/Y DFFSR_73/R DFFSR_23/S DFFSR_120/D INVX1_3/gnd DFFSR_23/S
+ DFFSR
XFILL_12_2 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_14_DFFSR_12 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_4_DFFSR_117 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_1_BUFX2_47 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_45_DFFSR_148 INVX1_67/gnd DFFSR_175/S FILL
XFILL_8_DFFSR_224 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_0_NAND3X1_11 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_35_DFFSR_151 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_8_DFFSR_5 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_49_DFFSR_255 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_9_OAI21X1_112 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_25_DFFSR_154 BUFX2_99/A DFFSR_7/S FILL
XFILL_39_DFFSR_258 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_49_DFFSR_29 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_38_DFFSR_69 BUFX2_98/A DFFSR_32/S FILL
XFILL_1_INVX1_201 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_7_NAND3X1_190 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_15_DFFSR_157 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_29_0_1 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_29_DFFSR_261 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_0_NAND3X1_1 BUFX2_98/A DFFSR_6/S FILL
XINVX1_13 INVX1_13/A DFFSR_4/gnd INVX1_13/Y DFFSR_98/S INVX1
XFILL_19_DFFSR_264 DFFSR_4/gnd DFFSR_98/S FILL
XDFFSR_66 DFFSR_66/Q DFFSR_82/CLK DFFSR_15/R DFFSR_5/S DFFSR_66/D BUFX2_77/gnd DFFSR_5/S
+ DFFSR
XFILL_0_NAND2X1_171 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_22_DFFSR_19 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_5_DFFSR_26 BUFX2_79/A DFFSR_6/S FILL
XFILL_11_DFFSR_59 AND2X2_38/B DFFSR_59/S FILL
XFILL_27_2_2 INVX1_3/gnd DFFSR_79/S FILL
XFILL_0_NOR2X1_36 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_6_OR2X2_5 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_9_1_1 XOR2X1_1/gnd DFFSR_208/S FILL
XINVX1_131 BUFX2_52/Y BUFX2_7/gnd INVX1_131/Y DFFSR_216/S INVX1
XFILL_8_NAND3X1_124 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_4_NOR2X1_7 BUFX2_98/A DFFSR_32/S FILL
XFILL_12_DFFPOSX1_28 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_1_DFFSR_154 BUFX2_99/A DFFSR_7/S FILL
XFILL_32_DFFSR_9 BUFX2_79/A DFFSR_6/S FILL
XFILL_1_NAND2X1_105 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_4_INVX1_128 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_42_DFFSR_185 INVX1_39/gnd DFFSR_54/S FILL
XFILL_46_DFFSR_76 BUFX2_79/A DFFSR_7/S FILL
XFILL_7_3_2 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_5_DFFSR_261 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_32_DFFSR_188 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_22_DFFSR_191 INVX1_67/gnd DFFSR_175/S FILL
XFILL_30_DFFSR_26 BUFX2_79/A DFFSR_6/S FILL
XFILL_2_INVX1_20 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_2_DFFSR_73 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_19_DFFSR_66 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_12_DFFSR_194 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_22_DFFPOSX1_17 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_1_BUFX2_11 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_6_NAND3X1_220 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_6_XOR2X1_3 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_54_5_0 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_45_DFFSR_112 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_2_DFFPOSX1_39 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_8_DFFSR_188 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_35_DFFSR_115 INVX1_1/gnd DFFSR_97/S FILL
XFILL_49_DFFSR_219 INVX1_67/gnd DFFSR_175/S FILL
XAND2X2_35 AND2X2_35/A AND2X2_35/B DFFSR_34/gnd AND2X2_35/Y DFFSR_34/S AND2X2
XFILL_25_DFFSR_118 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_39_DFFSR_222 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_38_DFFSR_33 BUFX2_98/A DFFSR_32/S FILL
XFILL_1_INVX1_165 BUFX2_99/A DFFSR_92/S FILL
XFILL_27_DFFSR_73 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_4_AND2X2_32 AND2X2_38/B DFFSR_23/S FILL
XFILL_7_NAND3X1_154 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_15_DFFSR_121 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_29_DFFSR_225 INVX1_67/gnd DFFSR_175/S FILL
XFILL_0_NAND2X1_135 DFFSR_34/gnd DFFSR_34/S FILL
XDFFSR_30 DFFSR_30/Q DFFSR_92/CLK DFFSR_2/R DFFSR_32/S DFFSR_6/Q BUFX2_98/A DFFSR_32/S
+ DFFSR
XFILL_19_DFFSR_228 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_11_DFFSR_23 AND2X2_38/B DFFSR_23/S FILL
XFILL_8_OAI22X1_8 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_2_NOR3X1_4 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_1_DFFSR_118 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_34_2 INVX1_1/gnd DFFSR_53/S FILL
XFILL_21_DFFPOSX1_47 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_42_DFFSR_149 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_46_DFFSR_40 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_35_DFFSR_80 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_5_DFFSR_225 INVX1_67/gnd DFFSR_175/S FILL
XFILL_32_DFFSR_152 INVX1_1/gnd DFFSR_53/S FILL
XFILL_46_DFFSR_256 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_22_DFFSR_155 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_2_DFFSR_37 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_36_DFFSR_259 BUFX2_79/A DFFSR_6/S FILL
XFILL_19_DFFSR_30 BUFX2_98/A DFFSR_32/S FILL
XFILL_6_BUFX2_65 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_12_DFFSR_158 INVX1_3/gnd DFFSR_23/S FILL
XFILL_26_DFFSR_262 BUFX2_98/A DFFSR_32/S FILL
XFILL_8_OAI21X1_106 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_16_DFFSR_265 INVX1_67/gnd DFFSR_175/S FILL
XFILL_20_CLKBUF1_20 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_6_NAND3X1_184 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_19_DFFSR_3 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_19_CLKBUF1_23 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_43_DFFSR_87 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_8_DFFSR_152 INVX1_1/gnd DFFSR_53/S FILL
XFILL_49_DFFSR_183 INVX1_67/gnd DFFSR_175/S FILL
XFILL_18_CLKBUF1_26 INVX1_1/gnd DFFSR_53/S FILL
XNAND3X1_220 NAND2X1_90/A NAND3X1_218/Y NAND3X1_219/Y DFFSR_46/gnd NAND2X1_99/B DFFSR_54/S
+ NAND3X1
XFILL_39_DFFSR_186 BUFX2_99/A DFFSR_92/S FILL
XFILL_17_CLKBUF1_29 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_27_DFFSR_37 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_1_INVX1_129 AND2X2_38/B DFFSR_23/S FILL
XFILL_16_DFFSR_77 BUFX2_98/A DFFSR_32/S FILL
XFILL_2_DFFSR_262 BUFX2_98/A DFFSR_32/S FILL
XFILL_7_NAND3X1_118 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_29_DFFSR_189 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_16_CLKBUF1_32 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_3_BUFX2_4 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_11_DFFPOSX1_22 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_15_CLKBUF1_35 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_19_DFFSR_192 INVX1_1/gnd DFFSR_97/S FILL
XNOR2X1_74 BUFX2_39/Y NOR2X1_74/B DFFSR_62/gnd NOR2X1_74/Y DFFSR_208/S NOR2X1
XFILL_14_CLKBUF1_38 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_13_CLKBUF1_41 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_4_NOR2X1_71 INVX1_1/gnd DFFSR_97/S FILL
XFILL_12_CLKBUF1_44 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_21_DFFPOSX1_11 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_42_DFFSR_113 BUFX2_99/A DFFSR_92/S FILL
XFILL_7_DFFSR_91 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_35_DFFSR_44 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_11_CLKBUF1_47 BUFX2_98/A DFFSR_32/S FILL
XFILL_24_DFFSR_84 BUFX2_99/A DFFSR_7/S FILL
XFILL_28_3_0 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_5_DFFSR_189 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_32_DFFSR_116 INVX1_3/gnd DFFSR_23/S FILL
XFILL_46_DFFSR_220 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_5_NAND3X1_214 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_22_DFFSR_119 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_36_DFFSR_223 INVX1_39/gnd DFFSR_34/S FILL
XFILL_1_DFFPOSX1_33 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_1_AND2X2_33 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_26_5_1 INVX1_3/gnd DFFSR_23/S FILL
XFILL_12_DFFSR_122 BUFX2_79/A DFFSR_7/S FILL
XFILL_6_BUFX2_29 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_26_DFFSR_226 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_2_AOI21X1_1 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_8_4_0 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_16_DFFSR_229 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_6_NAND3X1_148 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_6_6_1 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_32_DFFSR_91 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_8_DFFSR_116 INVX1_3/gnd DFFSR_23/S FILL
XFILL_43_DFFSR_51 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_5_OAI22X1_9 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_49_DFFSR_147 DFFSR_1/gnd DFFSR_1/S FILL
XNAND3X1_184 AOI21X1_27/C AOI21X1_27/B AOI21X1_27/A BUFX2_8/gnd AOI21X1_22/B DFFSR_51/S
+ NAND3X1
XFILL_39_DFFSR_150 AND2X2_38/B DFFSR_23/S FILL
XFILL_16_DFFSR_41 BUFX2_98/A DFFSR_6/S FILL
XFILL_2_DFFSR_226 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_29_DFFSR_153 INVX1_67/gnd DFFSR_201/S FILL
XFILL_3_BUFX2_76 OR2X2_2/gnd DFFSR_216/S FILL
XNAND3X1_3 BUFX2_82/A AND2X2_3/Y BUFX2_20/Y BUFX2_99/A AND2X2_6/A DFFSR_92/S NAND3X1
XFILL_43_DFFSR_257 INVX1_39/gnd DFFSR_34/S FILL
XFILL_20_DFFPOSX1_41 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_19_DFFSR_156 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_33_DFFSR_260 BUFX2_77/gnd DFFSR_5/S FILL
XNOR2X1_38 NOR2X1_38/A NOR2X1_38/B INVX1_3/gnd NOR2X1_38/Y DFFSR_79/S NOR2X1
XFILL_4_NAND3X1_244 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_23_DFFSR_263 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_40_DFFSR_98 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_4_NOR2X1_35 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_13_DFFSR_266 INVX1_67/gnd DFFSR_201/S FILL
XFILL_1_AND2X2_7 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_7_OAI21X1_100 INVX1_3/gnd DFFSR_79/S FILL
XFILL_7_DFFSR_55 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_24_DFFSR_48 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_13_DFFSR_88 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_11_CLKBUF1_11 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_5_DFFSR_153 INVX1_67/gnd DFFSR_201/S FILL
XFILL_36_0_1 BUFX2_99/A DFFSR_92/S FILL
XFILL_5_NAND3X1_178 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_46_DFFSR_184 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_10_CLKBUF1_14 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_9_DFFSR_260 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_36_DFFSR_187 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_34_2_2 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_9_CLKBUF1_17 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_26_DFFSR_190 INVX1_39/gnd DFFSR_34/S FILL
XFILL_7_DFFSR_2 BUFX2_79/A DFFSR_7/S FILL
XFILL_16_DFFSR_193 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_8_CLKBUF1_20 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_6_NAND3X1_112 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_7_CLKBUF1_23 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_10_DFFPOSX1_16 INVX1_67/gnd DFFSR_175/S FILL
XFILL_43_DFFSR_15 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_32_DFFSR_55 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_21_DFFSR_95 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_1_NOR2X1_72 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_6_CLKBUF1_26 INVX1_1/gnd DFFSR_53/S FILL
XFILL_49_DFFSR_111 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_5_CLKBUF1_29 XOR2X1_4/gnd DFFSR_91/S FILL
XNAND3X1_148 AOI21X1_14/A AOI21X1_14/B AOI21X1_8/Y BUFX2_8/gnd AOI21X1_15/B DFFSR_81/S
+ NAND3X1
XFILL_39_DFFSR_114 NOR3X1_6/gnd DFFSR_91/S FILL
XCLKBUF1_26 BUFX2_4/Y INVX1_1/gnd DFFSR_9/CLK DFFSR_53/S CLKBUF1
XFILL_4_CLKBUF1_32 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_5_OR2X2_2 OR2X2_2/gnd DFFSR_216/S FILL
XOR2X2_6 OR2X2_6/A OR2X2_6/B OR2X2_6/gnd OR2X2_6/Y DFFSR_53/S OR2X2
XFILL_2_DFFSR_190 INVX1_39/gnd DFFSR_34/S FILL
XFILL_29_DFFSR_117 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_3_BUFX2_40 INVX1_1/gnd DFFSR_97/S FILL
XFILL_43_DFFSR_221 AND2X2_38/B DFFSR_59/S FILL
XFILL_3_CLKBUF1_35 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_8_AND2X2_31 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_19_DFFSR_120 INVX1_3/gnd DFFSR_23/S FILL
XFILL_33_DFFSR_224 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_2_CLKBUF1_38 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_31_DFFSR_6 BUFX2_79/A DFFSR_6/S FILL
XFILL_23_DFFSR_227 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_1_CLKBUF1_41 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_4_NAND3X1_208 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_1_INVX1_96 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_40_DFFSR_62 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_13_DFFSR_230 INVX1_67/gnd DFFSR_201/S FILL
XFILL_0_CLKBUF1_44 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_0_DFFPOSX1_27 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_7_DFFSR_19 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_24_DFFSR_12 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_13_DFFSR_52 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_5_DFFSR_117 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_0_BUFX2_87 INVX1_1/gnd DFFSR_53/S FILL
XFILL_46_DFFSR_148 INVX1_67/gnd DFFSR_175/S FILL
XFILL_5_NAND3X1_142 INVX1_67/gnd DFFSR_175/S FILL
XFILL_9_DFFSR_224 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_36_DFFSR_151 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_50_DFFSR_255 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_26_DFFSR_154 BUFX2_99/A DFFSR_7/S FILL
XFILL_40_DFFSR_258 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_48_DFFSR_69 BUFX2_98/A DFFSR_32/S FILL
XFILL_2_INVX1_201 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_16_DFFSR_157 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_30_DFFSR_261 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_1_NAND3X1_1 BUFX2_98/A DFFSR_6/S FILL
XFILL_20_DFFSR_264 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_32_DFFSR_19 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_4_INVX1_13 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_4_DFFSR_66 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_10_DFFSR_99 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_21_DFFSR_59 AND2X2_38/B DFFSR_59/S FILL
XFILL_19_DFFPOSX1_35 INVX1_39/gnd DFFSR_54/S FILL
XFILL_1_NOR2X1_36 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_10_DFFSR_267 XOR2X1_1/gnd DFFSR_208/S FILL
XNAND3X1_112 NOR2X1_50/Y NOR2X1_51/Y NOR2X1_52/Y DFFSR_1/gnd XOR2X1_14/B DFFSR_1/S
+ NAND3X1
XFILL_3_NAND3X1_238 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_2_DFFSR_154 BUFX2_99/A DFFSR_7/S FILL
XFILL_43_DFFSR_185 INVX1_39/gnd DFFSR_54/S FILL
XFILL_6_DFFSR_261 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_33_DFFSR_188 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_23_DFFSR_191 INVX1_67/gnd DFFSR_175/S FILL
XFILL_4_NAND3X1_172 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_29_DFFSR_66 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_40_DFFSR_26 BUFX2_79/A DFFSR_6/S FILL
XFILL_1_INVX1_60 INVX1_39/gnd DFFSR_34/S FILL
XFILL_13_DFFSR_194 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_9_DFFPOSX1_46 INVX1_39/gnd DFFSR_34/S FILL
XFILL_13_DFFSR_16 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_0_BUFX2_51 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_46_DFFSR_112 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_5_NAND3X1_106 INVX1_3/gnd DFFSR_23/S FILL
XFILL_9_DFFSR_188 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_36_DFFSR_115 INVX1_1/gnd DFFSR_97/S FILL
XFILL_50_DFFSR_219 INVX1_67/gnd DFFSR_175/S FILL
XFILL_26_DFFSR_118 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_40_DFFSR_222 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_48_DFFSR_33 BUFX2_98/A DFFSR_32/S FILL
XFILL_2_INVX1_165 BUFX2_99/A DFFSR_92/S FILL
XFILL_37_DFFSR_73 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_5_AND2X2_32 AND2X2_38/B DFFSR_23/S FILL
XFILL_16_DFFSR_121 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_30_DFFSR_225 INVX1_67/gnd DFFSR_175/S FILL
XFILL_20_DFFSR_228 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_4_DFFSR_30 BUFX2_98/A DFFSR_32/S FILL
XFILL_10_DFFSR_63 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_21_DFFSR_23 AND2X2_38/B DFFSR_23/S FILL
XFILL_2_BUFX2_1 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_10_DFFSR_231 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_35_3_0 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_3_NAND3X1_202 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_9_OAI22X1_8 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_2_DFFSR_118 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_33_5_1 INVX1_1/gnd DFFSR_53/S FILL
XFILL_43_DFFSR_149 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_45_DFFSR_80 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_6_DFFSR_225 INVX1_67/gnd DFFSR_175/S FILL
XFILL_33_DFFSR_152 INVX1_1/gnd DFFSR_53/S FILL
XFILL_47_DFFSR_256 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_23_DFFSR_155 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_4_NAND3X1_136 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_18_DFFSR_70 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_1_INVX1_24 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_29_DFFSR_30 BUFX2_98/A DFFSR_32/S FILL
XFILL_1_DFFSR_77 BUFX2_98/A DFFSR_32/S FILL
XFILL_37_DFFSR_259 BUFX2_79/A DFFSR_6/S FILL
XFILL_13_DFFSR_158 INVX1_3/gnd DFFSR_23/S FILL
XFILL_9_DFFPOSX1_10 INVX1_67/gnd DFFSR_201/S FILL
XFILL_27_DFFSR_262 BUFX2_98/A DFFSR_32/S FILL
XFILL_6_NAND2X1_172 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_17_DFFSR_265 INVX1_67/gnd DFFSR_175/S FILL
XFILL_22_DFFPOSX1_2 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_0_BUFX2_15 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_21_DFFPOSX1_5 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_5_XOR2X1_7 BUFX2_98/A DFFSR_6/S FILL
XFILL_43_DFFSR_9 BUFX2_79/A DFFSR_6/S FILL
XFILL_9_DFFSR_152 INVX1_1/gnd DFFSR_53/S FILL
XFILL_18_DFFPOSX1_29 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_20_DFFPOSX1_8 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_50_DFFSR_183 INVX1_67/gnd DFFSR_175/S FILL
XFILL_40_DFFSR_186 BUFX2_99/A DFFSR_92/S FILL
XFILL_37_DFFSR_37 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_9_DFFSR_84 BUFX2_99/A DFFSR_7/S FILL
XFILL_2_INVX1_129 AND2X2_38/B DFFSR_23/S FILL
XFILL_26_DFFSR_77 BUFX2_98/A DFFSR_32/S FILL
XFILL_2_NAND3X1_232 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_3_DFFSR_262 BUFX2_98/A DFFSR_32/S FILL
XFILL_30_DFFSR_189 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_20_DFFSR_192 INVX1_1/gnd DFFSR_97/S FILL
XFILL_10_DFFSR_27 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_10_DFFSR_195 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_43_0_1 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_5_NOR2X1_71 INVX1_1/gnd DFFSR_97/S FILL
XFILL_3_NAND3X1_166 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_18_NOR3X1_1 INVX1_3/gnd DFFSR_79/S FILL
XFILL_43_DFFSR_113 BUFX2_99/A DFFSR_92/S FILL
XFILL_8_DFFPOSX1_40 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_45_DFFSR_44 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_41_2_2 BUFX2_98/A DFFSR_32/S FILL
XFILL_34_DFFSR_84 BUFX2_99/A DFFSR_7/S FILL
XFILL_6_DFFSR_189 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_33_DFFSR_116 INVX1_3/gnd DFFSR_23/S FILL
XFILL_47_DFFSR_220 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_23_DFFSR_119 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_4_NAND3X1_100 AND2X2_38/B DFFSR_59/S FILL
XFILL_1_DFFSR_41 BUFX2_98/A DFFSR_6/S FILL
XFILL_18_DFFSR_34 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_37_DFFSR_223 INVX1_39/gnd DFFSR_34/S FILL
XFILL_2_AND2X2_33 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_13_DFFSR_122 BUFX2_79/A DFFSR_7/S FILL
XFILL_5_BUFX2_69 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_27_DFFSR_226 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_3_AOI21X1_1 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_6_NAND2X1_136 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_17_DFFSR_229 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_11_XOR2X1_4 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_42_DFFSR_91 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_9_DFFSR_116 INVX1_3/gnd DFFSR_23/S FILL
XNAND2X1_172 NAND3X1_8/Y NAND3X1_72/Y OR2X2_1/gnd INVX1_211/A DFFSR_59/S NAND2X1
XFILL_6_OAI22X1_9 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_4_OAI21X1_118 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_50_DFFSR_147 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_8_AOI21X1_64 AND2X2_38/B DFFSR_59/S FILL
XFILL_27_DFFPOSX1_48 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_40_DFFSR_150 AND2X2_38/B DFFSR_23/S FILL
XFILL_9_DFFSR_48 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_7_AOI21X1_67 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_26_DFFSR_41 BUFX2_98/A DFFSR_6/S FILL
XFILL_15_DFFSR_81 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_2_NAND3X1_196 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_3_DFFSR_226 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_30_DFFSR_153 INVX1_67/gnd DFFSR_201/S FILL
XFILL_6_AOI21X1_70 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_44_DFFSR_257 INVX1_39/gnd DFFSR_34/S FILL
XFILL_20_DFFSR_156 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_34_DFFSR_260 BUFX2_77/gnd DFFSR_5/S FILL
XAOI21X1_70 OR2X2_6/Y XOR2X1_15/Y AOI21X1_70/C OR2X2_6/gnd AOI21X1_70/Y DFFSR_92/S
+ AOI21X1
XFILL_10_DFFSR_159 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_24_DFFSR_263 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_50_DFFSR_98 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_5_NOR2X1_35 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_3_NAND3X1_130 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_14_DFFSR_266 INVX1_67/gnd DFFSR_201/S FILL
XFILL_30_DFFSR_3 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_34_DFFSR_48 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_23_DFFSR_88 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_6_DFFSR_95 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_5_NAND2X1_166 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_6_DFFSR_153 INVX1_67/gnd DFFSR_201/S FILL
XFILL_47_DFFSR_184 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_37_DFFSR_187 DFFSR_1/gnd DFFSR_81/S FILL
XBUFX2_73 BUFX2_73/A OR2X2_6/gnd dout[2] DFFSR_92/S BUFX2
XFILL_5_BUFX2_33 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_0_DFFSR_263 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_10_DFFPOSX1_2 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_17_DFFPOSX1_23 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_27_DFFSR_190 INVX1_39/gnd DFFSR_34/S FILL
XFILL_6_NAND2X1_100 INVX1_39/gnd DFFSR_54/S FILL
XFILL_17_DFFSR_193 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_1_NAND3X1_226 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_9_DFFPOSX1_5 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_42_DFFSR_55 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_3_INVX1_89 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_31_DFFSR_95 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_8_DFFPOSX1_8 OR2X2_4/gnd DFFSR_32/S FILL
XNAND2X1_136 DFFSR_276/S INVX1_194/A BUFX2_72/gnd NAND2X1_136/Y DFFSR_276/S NAND2X1
XFILL_2_NOR2X1_72 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_50_DFFSR_111 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_8_AOI21X1_28 AND2X2_38/B DFFSR_23/S FILL
XFILL_27_DFFPOSX1_12 AND2X2_38/B DFFSR_23/S FILL
XFILL_40_DFFSR_114 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_9_DFFSR_12 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_7_AOI21X1_31 INVX1_39/gnd DFFSR_34/S FILL
XFILL_15_DFFSR_45 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_2_NAND3X1_160 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_3_DFFSR_190 INVX1_39/gnd DFFSR_34/S FILL
XFILL_30_DFFSR_117 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_2_BUFX2_80 BUFX2_79/A DFFSR_6/S FILL
XFILL_15_0_2 INVX1_39/gnd DFFSR_34/S FILL
XFILL_44_DFFSR_221 AND2X2_38/B DFFSR_59/S FILL
XFILL_6_AOI21X1_34 INVX1_39/gnd DFFSR_34/S FILL
XFILL_9_AND2X2_31 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_7_DFFPOSX1_34 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_20_DFFSR_120 INVX1_3/gnd DFFSR_23/S FILL
XFILL_5_AOI21X1_37 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_34_DFFSR_224 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_10_DFFSR_123 XOR2X1_4/gnd DFFSR_97/S FILL
XAOI21X1_34 AOI21X1_34/A AOI21X1_41/B OAI21X1_74/Y INVX1_39/gnd OAI22X1_51/C DFFSR_34/S
+ AOI21X1
XFILL_4_AOI21X1_40 INVX1_39/gnd DFFSR_54/S FILL
XFILL_24_DFFSR_227 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_0_AOI21X1_2 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_50_DFFSR_62 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_3_AOI21X1_43 INVX1_3/gnd DFFSR_79/S FILL
XFILL_14_DFFSR_230 INVX1_67/gnd DFFSR_201/S FILL
XFILL_2_AOI21X1_46 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_34_DFFSR_12 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_23_DFFSR_52 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_6_DFFSR_59 AND2X2_38/B DFFSR_59/S FILL
XFILL_5_NAND2X1_130 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_1_AOI21X1_49 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_6_DFFSR_117 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_12_DFFSR_92 BUFX2_99/A DFFSR_92/S FILL
XFILL_47_DFFSR_148 INVX1_67/gnd DFFSR_175/S FILL
XFILL_0_AOI21X1_52 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_37_DFFSR_151 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_0_DFFSR_227 BUFX2_7/gnd DFFSR_151/S FILL
XBUFX2_37 rst INVX1_1/gnd NOR3X1_6/A DFFSR_97/S BUFX2
XFILL_27_DFFSR_154 BUFX2_99/A DFFSR_7/S FILL
XFILL_3_OAI21X1_112 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_26_DFFPOSX1_42 INVX1_39/gnd DFFSR_34/S FILL
XFILL_41_DFFSR_258 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_42_3_0 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_3_INVX1_201 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_17_DFFSR_157 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_8_OAI21X1_76 INVX1_1/gnd DFFSR_53/S FILL
XFILL_1_NAND3X1_190 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_31_DFFSR_261 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_2_NAND3X1_1 BUFX2_98/A DFFSR_6/S FILL
XFILL_6_NAND2X1_97 INVX1_1/gnd DFFSR_97/S FILL
XFILL_7_OAI21X1_79 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_21_DFFSR_264 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_42_DFFSR_19 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_3_INVX1_53 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_40_5_1 BUFX2_98/A DFFSR_6/S FILL
XFILL_20_DFFSR_99 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_31_DFFSR_59 AND2X2_38/B DFFSR_59/S FILL
XFILL_2_NOR2X1_36 OR2X2_1/gnd DFFSR_51/S FILL
XNAND2X1_100 AOI21X1_34/A AOI21X1_41/B INVX1_39/gnd OAI21X1_75/B DFFSR_54/S NAND2X1
XFILL_6_OAI21X1_82 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_11_DFFSR_267 XOR2X1_1/gnd DFFSR_208/S FILL
XNAND2X1_97 INVX1_135/A AOI22X1_25/B INVX1_1/gnd NOR2X1_71/B DFFSR_97/S NAND2X1
XFILL_5_OAI21X1_85 INVX1_39/gnd DFFSR_54/S FILL
XOAI21X1_82 OAI21X1_82/A AOI21X1_38/Y INVX1_171/Y DFFSR_28/gnd AOI21X1_45/A DFFSR_8/S
+ OAI21X1
XFILL_2_NAND3X1_124 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_4_OAI21X1_88 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_3_DFFSR_154 BUFX2_99/A DFFSR_7/S FILL
XFILL_2_BUFX2_44 INVX1_3/gnd DFFSR_79/S FILL
XFILL_44_DFFSR_185 INVX1_39/gnd DFFSR_54/S FILL
XFILL_3_OAI21X1_91 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_7_DFFSR_261 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_4_NAND2X1_160 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_34_DFFSR_188 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_2_OAI21X1_94 INVX1_67/gnd DFFSR_175/S FILL
XFILL_24_DFFSR_191 INVX1_67/gnd DFFSR_175/S FILL
XFILL_1_OAI21X1_97 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_39_DFFSR_66 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_50_DFFSR_26 BUFX2_79/A DFFSR_6/S FILL
XFILL_14_DFFSR_194 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_16_DFFPOSX1_17 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_2_AOI21X1_10 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_23_DFFSR_16 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_6_DFFSR_23 AND2X2_38/B DFFSR_23/S FILL
XFILL_12_DFFSR_56 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_1_AOI21X1_13 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_47_DFFSR_112 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_0_NAND3X1_220 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_0_AOI21X1_16 INVX1_67/gnd DFFSR_175/S FILL
XFILL_37_DFFSR_115 INVX1_1/gnd DFFSR_97/S FILL
XFILL_5_NOR2X1_4 INVX1_1/gnd DFFSR_53/S FILL
XFILL_0_DFFSR_191 INVX1_67/gnd DFFSR_175/S FILL
XFILL_27_DFFSR_118 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_42_DFFSR_6 BUFX2_79/A DFFSR_6/S FILL
XFILL_9_OAI21X1_37 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_41_DFFSR_222 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_3_INVX1_165 BUFX2_99/A DFFSR_92/S FILL
XFILL_6_AND2X2_32 AND2X2_38/B DFFSR_23/S FILL
XFILL_47_DFFSR_73 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_17_DFFSR_121 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_50_0_1 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_8_OAI21X1_40 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_31_DFFSR_225 INVX1_67/gnd DFFSR_175/S FILL
XFILL_1_NAND3X1_154 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_6_NAND2X1_61 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_7_OAI21X1_43 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_21_DFFSR_228 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_3_DFFSR_70 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_3_INVX1_17 AND2X2_38/B DFFSR_59/S FILL
XFILL_20_DFFSR_63 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_31_DFFSR_23 AND2X2_38/B DFFSR_23/S FILL
XFILL_6_DFFPOSX1_28 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_48_2_2 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_6_OAI21X1_46 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_5_NAND2X1_64 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_11_DFFSR_231 DFFSR_46/gnd DFFSR_62/S FILL
XNAND2X1_61 OR2X2_2/B OR2X2_2/A OR2X2_2/gnd OAI21X1_26/C DFFSR_216/S NAND2X1
XFILL_4_NAND2X1_67 AND2X2_38/B DFFSR_59/S FILL
XFILL_5_OAI21X1_49 DFFSR_34/gnd DFFSR_1/S FILL
XOAI21X1_46 INVX1_152/A OAI21X1_41/A OAI21X1_46/C DFFSR_34/gnd OAI21X1_54/C DFFSR_1/S
+ OAI21X1
XFILL_3_NAND2X1_70 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_3_DFFSR_118 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_4_OAI21X1_52 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_44_DFFSR_149 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_15_DFFPOSX1_47 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_2_NAND2X1_73 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_3_OAI21X1_55 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_7_DFFSR_225 INVX1_67/gnd DFFSR_175/S FILL
XFILL_4_NAND2X1_124 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_34_DFFSR_152 INVX1_1/gnd DFFSR_53/S FILL
XFILL_48_DFFSR_256 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_1_NAND2X1_76 INVX1_3/gnd DFFSR_23/S FILL
XFILL_2_OAI21X1_58 INVX1_39/gnd DFFSR_54/S FILL
XFILL_11_AOI22X1_24 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_55_10 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_24_DFFSR_155 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_1_OAI21X1_61 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_0_NAND2X1_79 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_0_INVX1_202 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_28_DFFSR_70 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_39_DFFSR_30 BUFX2_98/A DFFSR_32/S FILL
XFILL_38_DFFSR_259 BUFX2_79/A DFFSR_6/S FILL
XFILL_10_AOI22X1_27 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_0_INVX1_64 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_14_DFFSR_158 INVX1_3/gnd DFFSR_23/S FILL
XFILL_0_OAI21X1_64 INVX1_1/gnd DFFSR_53/S FILL
XFILL_16_1_0 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_28_DFFSR_262 BUFX2_98/A DFFSR_32/S FILL
XFILL_2_OAI21X1_106 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_18_DFFSR_265 INVX1_67/gnd DFFSR_175/S FILL
XFILL_25_DFFPOSX1_36 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_12_DFFSR_20 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_14_3_1 INVX1_39/gnd DFFSR_54/S FILL
XFILL_0_NAND3X1_184 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_9_NAND3X1_239 DFFSR_8/gnd DFFSR_60/S FILL
XNOR2X1_8 NOR2X1_8/A NOR2X1_8/B OR2X2_6/gnd NOR2X1_8/Y DFFSR_92/S NOR2X1
XFILL_3_NOR3X1_1 INVX1_3/gnd DFFSR_79/S FILL
XDFFSR_265 DFFSR_265/Q CLKBUF1_47/Y DFFSR_266/R DFFSR_175/S DFFSR_265/D INVX1_67/gnd
+ DFFSR_175/S DFFSR
XFILL_0_DFFSR_155 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_12_5_2 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_41_DFFSR_186 BUFX2_99/A DFFSR_92/S FILL
XFILL_3_INVX1_129 AND2X2_38/B DFFSR_23/S FILL
XFILL_47_DFFSR_37 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_36_DFFSR_77 BUFX2_98/A DFFSR_32/S FILL
XFILL_4_DFFSR_262 BUFX2_98/A DFFSR_32/S FILL
XFILL_31_DFFSR_189 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_1_NAND3X1_118 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_6_NAND2X1_25 BUFX2_99/A DFFSR_7/S FILL
XFILL_21_DFFSR_192 INVX1_1/gnd DFFSR_97/S FILL
XFILL_3_DFFSR_34 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_20_DFFSR_27 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_3_NAND2X1_154 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_6_OAI21X1_10 BUFX2_79/A DFFSR_7/S FILL
XFILL_5_NAND2X1_28 AND2X2_38/B DFFSR_59/S FILL
XFILL_11_DFFSR_195 DFFSR_46/gnd DFFSR_62/S FILL
XNAND2X1_25 DFFSR_120/D NOR2X1_5/Y BUFX2_99/A OAI21X1_8/C DFFSR_7/S NAND2X1
XFILL_4_NAND2X1_31 INVX1_3/gnd DFFSR_23/S FILL
XFILL_5_OAI21X1_13 INVX1_39/gnd DFFSR_54/S FILL
XFILL_6_NOR2X1_71 INVX1_1/gnd DFFSR_97/S FILL
XFILL_8_5 BUFX2_7/gnd DFFSR_151/S FILL
XOAI21X1_10 INVX1_75/Y OAI21X1_9/B OAI21X1_10/C BUFX2_79/A NOR2X1_39/B DFFSR_7/S OAI21X1
XFILL_4_OAI21X1_16 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_3_NAND2X1_34 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_9_DFFSR_9 BUFX2_79/A DFFSR_6/S FILL
XDFFPOSX1_28 DFFPOSX1_28/Q CLKBUF1_43/Y AOI21X1_50/Y BUFX2_72/gnd DFFSR_201/S DFFPOSX1
XFILL_44_DFFSR_113 BUFX2_99/A DFFSR_92/S FILL
XFILL_2_NAND2X1_37 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_15_DFFPOSX1_11 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_3_OAI21X1_19 BUFX2_98/A DFFSR_32/S FILL
XFILL_44_DFFSR_84 BUFX2_99/A DFFSR_7/S FILL
XFILL_7_DFFSR_189 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_34_DFFSR_116 INVX1_3/gnd DFFSR_23/S FILL
XFILL_9_NAND3X1_93 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_48_DFFSR_220 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_1_NAND2X1_40 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_2_OAI21X1_22 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_24_DFFSR_119 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_8_NAND3X1_96 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_0_NAND2X1_43 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_1_OAI21X1_25 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_0_INVX1_28 DFFSR_28/gnd DFFSR_3/S FILL
XAOI21X1_4 NOR3X1_4/B NOR3X1_4/A BUFX2_40/Y BUFX2_98/A AOI21X1_4/Y DFFSR_32/S AOI21X1
XFILL_0_INVX1_166 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_0_DFFSR_81 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_28_DFFSR_34 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_38_DFFSR_223 INVX1_39/gnd DFFSR_34/S FILL
XFILL_17_DFFSR_74 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_3_AND2X2_33 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_14_DFFSR_122 BUFX2_79/A DFFSR_7/S FILL
XFILL_7_NAND3X1_99 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_0_OAI21X1_28 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_28_DFFSR_226 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_4_AOI21X1_1 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_18_DFFSR_229 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_0_NAND3X1_148 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_22_0_2 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_7_OAI22X1_9 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_5_DFFPOSX1_22 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_0_DFFSR_119 OR2X2_4/gnd DFFSR_3/S FILL
XDFFSR_229 DFFSR_237/D CLKBUF1_12/Y BUFX2_70/Y DFFSR_59/S DFFSR_229/D OR2X2_1/gnd
+ DFFSR_59/S DFFSR
XFILL_30_6 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_41_DFFSR_150 AND2X2_38/B DFFSR_23/S FILL
XFILL_8_DFFSR_88 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_36_DFFSR_41 BUFX2_98/A DFFSR_6/S FILL
XFILL_25_DFFSR_81 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_47_1 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_4_DFFSR_226 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_31_DFFSR_153 INVX1_67/gnd DFFSR_201/S FILL
XFILL_2_1_2 INVX1_67/gnd DFFSR_201/S FILL
XFILL_45_DFFSR_257 INVX1_39/gnd DFFSR_34/S FILL
XFILL_21_DFFSR_156 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_14_DFFPOSX1_41 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_35_DFFSR_260 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_3_AOI22X1_12 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_3_NAND2X1_118 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_11_DFFSR_159 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_25_DFFSR_263 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_2_AOI22X1_15 DFFSR_46/gnd DFFSR_54/S FILL
XINVX1_2 INVX1_2/A OR2X2_6/gnd INVX1_2/Y DFFSR_92/S INVX1
XFILL_6_NOR2X1_35 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_15_DFFSR_266 INVX1_67/gnd DFFSR_201/S FILL
XFILL_11_OAI22X1_36 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_1_AOI22X1_18 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_17_NOR3X1_5 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_10_OAI22X1_39 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_0_AOI22X1_21 AND2X2_38/B DFFSR_59/S FILL
XFILL_44_DFFSR_48 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_1_OAI21X1_100 INVX1_3/gnd DFFSR_79/S FILL
XFILL_7_DFFSR_153 INVX1_67/gnd DFFSR_201/S FILL
XFILL_33_DFFSR_88 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_49_3_0 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_24_DFFPOSX1_30 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_9_NAND3X1_57 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_48_DFFSR_184 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_8_NAND3X1_60 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_9_OAI22X1_42 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_0_DFFSR_45 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_8_NAND3X1_233 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_0_INVX1_130 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_38_DFFSR_187 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_17_DFFSR_38 BUFX2_98/A DFFSR_6/S FILL
XFILL_8_OAI22X1_45 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_7_NAND3X1_63 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_47_5_1 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_1_DFFSR_263 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_4_BUFX2_73 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_28_DFFSR_190 INVX1_39/gnd DFFSR_34/S FILL
XFILL_6_NAND3X1_66 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_7_OAI22X1_48 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_18_DFFSR_193 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_5_NAND3X1_69 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_6_OAI22X1_51 INVX1_39/gnd DFFSR_54/S FILL
XFILL_0_NAND3X1_112 DFFSR_1/gnd DFFSR_1/S FILL
XNAND3X1_66 DFFSR_153/D AND2X2_18/B BUFX2_27/Y BUFX2_7/gnd AND2X2_19/B DFFSR_151/S
+ NAND3X1
XFILL_10_XOR2X1_8 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_4_NAND3X1_72 INVX1_39/gnd DFFSR_34/S FILL
XFILL_41_DFFSR_95 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_3_NOR2X1_72 DFFSR_8/gnd DFFSR_60/S FILL
XOAI22X1_51 INVX1_131/Y NAND2X1_99/Y OAI22X1_51/C OAI22X1_51/D INVX1_39/gnd OAI22X1_51/Y
+ DFFSR_54/S OAI22X1
XFILL_51_DFFSR_111 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_3_NAND3X1_75 BUFX2_79/A DFFSR_7/S FILL
XDFFSR_193 DFFSR_201/D CLKBUF1_34/Y BUFX2_62/Y DFFSR_175/S DFFSR_193/D OR2X2_2/gnd
+ DFFSR_175/S DFFSR
XFILL_2_NAND2X1_148 INVX1_67/gnd DFFSR_175/S FILL
XFILL_2_AND2X2_4 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_41_DFFSR_114 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_8_DFFSR_52 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_2_NAND3X1_78 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_14_DFFSR_85 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_25_DFFSR_45 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_4_DFFSR_190 INVX1_39/gnd DFFSR_34/S FILL
XFILL_31_DFFSR_117 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_1_NAND3X1_81 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_45_DFFSR_221 AND2X2_38/B DFFSR_59/S FILL
XFILL_21_DFFSR_120 INVX1_3/gnd DFFSR_23/S FILL
XFILL_0_NAND3X1_84 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_35_DFFSR_224 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_0_AND2X2_34 AND2X2_38/B DFFSR_59/S FILL
XFILL_11_DFFSR_123 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_13_6_0 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_25_DFFSR_227 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_1_AOI21X1_2 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_15_DFFSR_230 INVX1_67/gnd DFFSR_201/S FILL
XFILL_20_DFFSR_7 BUFX2_79/A DFFSR_7/S FILL
XINVX1_86 INVX1_86/A DFFSR_46/gnd INVX1_86/Y DFFSR_54/S INVX1
XFILL_44_DFFSR_12 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_33_DFFSR_52 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_5_DFFSR_99 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_7_DFFSR_117 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_22_DFFSR_92 BUFX2_99/A DFFSR_92/S FILL
XFILL_48_DFFSR_148 INVX1_67/gnd DFFSR_175/S FILL
XFILL_8_NAND3X1_24 INVX1_1/gnd DFFSR_97/S FILL
XFILL_4_BUFX2_8 BUFX2_8/gnd DFFSR_51/S FILL
XINVX1_204 BUFX2_76/A BUFX2_7/gnd INVX1_204/Y DFFSR_216/S INVX1
XFILL_38_DFFSR_151 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_8_NAND3X1_197 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_1_DFFSR_227 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_7_NAND3X1_27 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_4_BUFX2_37 INVX1_1/gnd DFFSR_97/S FILL
XFILL_4_DFFPOSX1_16 INVX1_67/gnd DFFSR_175/S FILL
XFILL_28_DFFSR_154 BUFX2_99/A DFFSR_7/S FILL
XFILL_1_NAND2X1_178 INVX1_1/gnd DFFSR_53/S FILL
XFILL_42_DFFSR_258 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_4_INVX1_201 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_7_OAI22X1_12 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_6_NAND3X1_30 BUFX2_79/A DFFSR_6/S FILL
XFILL_18_DFFSR_157 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_32_DFFSR_261 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_6_OAI22X1_15 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_5_NAND3X1_33 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_41_DFFSR_3 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_3_NAND3X1_1 BUFX2_98/A DFFSR_6/S FILL
XNAND3X1_30 DFFSR_76/D BUFX2_18/Y NOR2X1_2/Y BUFX2_79/A NAND3X1_31/B DFFSR_6/S NAND3X1
XFILL_22_DFFSR_264 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_5_OAI22X1_18 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_4_NAND3X1_36 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_30_DFFSR_99 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_2_INVX1_93 INVX1_3/gnd DFFSR_23/S FILL
XFILL_41_DFFSR_59 AND2X2_38/B DFFSR_59/S FILL
XFILL_3_NOR2X1_36 OR2X2_1/gnd DFFSR_51/S FILL
XOAI22X1_15 INVX1_35/Y OAI22X1_6/B INVX1_36/Y OAI22X1_6/D DFFSR_28/gnd NOR2X1_19/A
+ DFFSR_3/S OAI22X1
XFILL_13_DFFPOSX1_35 INVX1_39/gnd DFFSR_54/S FILL
XFILL_3_NAND3X1_39 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_12_DFFSR_267 XOR2X1_1/gnd DFFSR_208/S FILL
XDFFSR_157 INVX1_95/A CLKBUF1_14/Y BUFX2_66/Y DFFSR_151/S DFFSR_157/D XOR2X1_1/gnd
+ DFFSR_151/S DFFSR
XFILL_4_OAI22X1_21 BUFX2_98/A DFFSR_32/S FILL
XFILL_2_NAND2X1_112 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_8_DFFSR_16 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_3_OAI22X1_24 BUFX2_98/A DFFSR_32/S FILL
XFILL_2_NAND3X1_42 BUFX2_79/A DFFSR_6/S FILL
XFILL_14_DFFSR_49 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_4_DFFSR_154 BUFX2_99/A DFFSR_7/S FILL
XFILL_2_OAI22X1_27 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_1_NAND3X1_45 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_1_BUFX2_84 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_45_DFFSR_185 INVX1_39/gnd DFFSR_54/S FILL
XFILL_23_1_0 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_0_NAND3X1_48 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_8_DFFSR_261 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_1_OAI22X1_30 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_35_DFFSR_188 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_23_DFFPOSX1_24 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_0_OAI22X1_33 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_25_DFFSR_191 INVX1_67/gnd DFFSR_175/S FILL
XFILL_21_3_1 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_49_DFFSR_66 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_15_DFFSR_194 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_7_NAND3X1_227 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_3_2_0 INVX1_67/gnd DFFSR_175/S FILL
XFILL_3_DFFPOSX1_46 INVX1_39/gnd DFFSR_34/S FILL
XINVX1_50 DFFSR_23/D BUFX2_98/A INVX1_50/Y DFFSR_6/S INVX1
XFILL_19_5_2 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_33_DFFSR_16 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_5_DFFSR_63 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_22_DFFSR_56 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_11_DFFSR_96 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_0_NOR2X1_73 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_48_DFFSR_112 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_1_4_1 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_38_DFFSR_115 INVX1_1/gnd DFFSR_97/S FILL
XINVX1_168 INVX1_168/A OR2X2_6/gnd INVX1_168/Y DFFSR_92/S INVX1
XFILL_8_NAND3X1_161 AND2X2_38/B DFFSR_23/S FILL
XFILL_1_DFFSR_191 INVX1_67/gnd DFFSR_175/S FILL
XFILL_28_DFFSR_118 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_1_NAND2X1_142 INVX1_67/gnd DFFSR_175/S FILL
XFILL_42_DFFSR_222 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_4_INVX1_165 BUFX2_99/A DFFSR_92/S FILL
XFILL_7_AND2X2_32 AND2X2_38/B DFFSR_23/S FILL
XFILL_18_DFFSR_121 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_32_DFFSR_225 INVX1_67/gnd DFFSR_175/S FILL
XFILL_22_DFFSR_228 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_30_DFFSR_63 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_2_INVX1_57 BUFX2_98/A DFFSR_32/S FILL
XFILL_41_DFFSR_23 AND2X2_38/B DFFSR_23/S FILL
XFILL_12_DFFSR_231 DFFSR_46/gnd DFFSR_62/S FILL
XDFFSR_121 BUFX2_82/A CLKBUF1_40/Y BUFX2_49/Y DFFSR_53/S INVX1_9/A OR2X2_6/gnd DFFSR_53/S
+ DFFSR
XFILL_12_3 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_14_DFFSR_13 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_4_DFFSR_118 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_1_BUFX2_48 AND2X2_38/B DFFSR_59/S FILL
XFILL_45_DFFSR_149 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_8_DFFSR_225 INVX1_67/gnd DFFSR_175/S FILL
XFILL_0_NAND3X1_12 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_8_DFFSR_6 BUFX2_79/A DFFSR_6/S FILL
XFILL_35_DFFSR_152 INVX1_1/gnd DFFSR_53/S FILL
XFILL_49_DFFSR_256 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_25_DFFSR_155 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_1_INVX1_202 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_49_DFFSR_30 BUFX2_98/A DFFSR_32/S FILL
XFILL_39_DFFSR_259 BUFX2_79/A DFFSR_6/S FILL
XFILL_38_DFFSR_70 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_29_0_2 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_15_DFFSR_158 INVX1_3/gnd DFFSR_23/S FILL
XFILL_7_NAND3X1_191 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_29_DFFSR_262 BUFX2_98/A DFFSR_32/S FILL
XFILL_0_NAND3X1_2 BUFX2_99/A DFFSR_7/S FILL
XFILL_3_DFFPOSX1_10 INVX1_67/gnd DFFSR_201/S FILL
XFILL_19_DFFSR_265 INVX1_67/gnd DFFSR_175/S FILL
XINVX1_14 DFFSR_34/D BUFX2_98/A INVX1_14/Y DFFSR_6/S INVX1
XFILL_0_NAND2X1_172 OR2X2_1/gnd DFFSR_59/S FILL
XDFFSR_67 DFFSR_67/Q DFFSR_1/CLK DFFSR_1/R DFFSR_34/S DFFSR_67/D DFFSR_34/gnd DFFSR_34/S
+ DFFSR
XFILL_5_DFFSR_27 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_11_DFFSR_60 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_22_DFFSR_20 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_0_NOR2X1_37 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_6_OR2X2_6 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_9_1_2 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_8_NAND3X1_125 BUFX2_77/gnd DFFSR_98/S FILL
XINVX1_132 BUFX2_57/Y NOR3X1_6/gnd INVX1_132/Y DFFSR_91/S INVX1
XFILL_4_NOR2X1_8 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_1_DFFSR_155 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_12_DFFPOSX1_29 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_1_NAND2X1_106 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_42_DFFSR_186 BUFX2_99/A DFFSR_92/S FILL
XFILL_46_DFFSR_77 BUFX2_98/A DFFSR_32/S FILL
XFILL_5_DFFSR_262 BUFX2_98/A DFFSR_32/S FILL
XFILL_32_DFFSR_189 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_22_DFFSR_192 INVX1_1/gnd DFFSR_97/S FILL
XFILL_30_DFFSR_27 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_2_DFFSR_74 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_2_INVX1_21 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_19_DFFSR_67 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_12_DFFSR_195 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_22_DFFPOSX1_18 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_1_BUFX2_12 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_6_NAND3X1_221 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_54_5_1 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_45_DFFSR_113 BUFX2_99/A DFFSR_92/S FILL
XFILL_6_XOR2X1_4 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_2_DFFPOSX1_40 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_8_DFFSR_189 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_35_DFFSR_116 INVX1_3/gnd DFFSR_23/S FILL
XAND2X2_36 INVX1_145/A INVX1_159/A NOR3X1_6/gnd AND2X2_36/Y DFFSR_79/S AND2X2
XFILL_49_DFFSR_220 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_25_DFFSR_119 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_1_INVX1_166 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_39_DFFSR_223 INVX1_39/gnd DFFSR_34/S FILL
XFILL_27_DFFSR_74 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_4_AND2X2_33 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_38_DFFSR_34 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_15_DFFSR_122 BUFX2_79/A DFFSR_7/S FILL
XFILL_7_NAND3X1_155 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_29_DFFSR_226 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_5_AOI21X1_1 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_0_NAND2X1_136 BUFX2_72/gnd DFFSR_276/S FILL
XDFFSR_31 DFFSR_23/D DFFSR_7/CLK DFFSR_9/R DFFSR_6/S DFFSR_7/Q BUFX2_79/A DFFSR_6/S
+ DFFSR
XFILL_19_DFFSR_229 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_11_DFFSR_24 BUFX2_98/A DFFSR_6/S FILL
XFILL_8_OAI22X1_9 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_2_NOR3X1_5 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_1_DFFSR_119 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_34_3 INVX1_1/gnd DFFSR_53/S FILL
XFILL_21_DFFPOSX1_48 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_20_6_0 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_42_DFFSR_150 AND2X2_38/B DFFSR_23/S FILL
XFILL_46_DFFSR_41 BUFX2_98/A DFFSR_6/S FILL
XFILL_35_DFFSR_81 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_5_DFFSR_226 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_32_DFFSR_153 INVX1_67/gnd DFFSR_201/S FILL
XFILL_46_DFFSR_257 INVX1_39/gnd DFFSR_34/S FILL
XFILL_22_DFFSR_156 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_36_DFFSR_260 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_2_DFFSR_38 BUFX2_98/A DFFSR_6/S FILL
XFILL_19_DFFSR_31 BUFX2_79/A DFFSR_6/S FILL
XFILL_12_DFFSR_159 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_6_BUFX2_66 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_26_DFFSR_263 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_8_OAI21X1_107 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_16_DFFSR_266 INVX1_67/gnd DFFSR_201/S FILL
XFILL_6_NAND3X1_185 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_20_CLKBUF1_21 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_12_XOR2X1_1 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_19_DFFSR_4 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_19_CLKBUF1_24 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_8_DFFSR_153 INVX1_67/gnd DFFSR_201/S FILL
XFILL_43_DFFSR_88 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_49_DFFSR_184 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_18_CLKBUF1_27 INVX1_1/gnd DFFSR_97/S FILL
XNAND3X1_221 INVX1_169/A NAND2X1_99/A NAND2X1_99/B DFFSR_46/gnd AOI21X1_34/A DFFSR_54/S
+ NAND3X1
XFILL_17_CLKBUF1_30 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_1_INVX1_130 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_39_DFFSR_187 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_16_DFFSR_78 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_27_DFFSR_38 BUFX2_98/A DFFSR_6/S FILL
XFILL_7_NAND3X1_119 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_2_DFFSR_263 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_16_CLKBUF1_33 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_29_DFFSR_190 INVX1_39/gnd DFFSR_34/S FILL
XFILL_11_DFFPOSX1_23 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_3_BUFX2_5 AND2X2_38/B DFFSR_59/S FILL
XFILL_19_DFFSR_193 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_15_CLKBUF1_36 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_0_NAND2X1_100 INVX1_39/gnd DFFSR_54/S FILL
XNOR2X1_75 BUFX2_8/Y BUFX2_35/Y BUFX2_8/gnd NOR2X1_75/Y DFFSR_51/S NOR2X1
XFILL_14_CLKBUF1_39 INVX1_1/gnd DFFSR_53/S FILL
XFILL_51_DFFSR_95 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_4_NOR2X1_72 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_13_CLKBUF1_42 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_30_1_0 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_12_CLKBUF1_45 BUFX2_79/A DFFSR_7/S FILL
XFILL_21_DFFPOSX1_12 AND2X2_38/B DFFSR_23/S FILL
XFILL_42_DFFSR_114 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_35_DFFSR_45 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_7_DFFSR_92 BUFX2_99/A DFFSR_92/S FILL
XFILL_11_CLKBUF1_48 INVX1_3/gnd DFFSR_79/S FILL
XFILL_24_DFFSR_85 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_28_3_1 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_5_DFFSR_190 INVX1_39/gnd DFFSR_34/S FILL
XFILL_32_DFFSR_117 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_46_DFFSR_221 AND2X2_38/B DFFSR_59/S FILL
XFILL_5_NAND3X1_215 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_22_DFFSR_120 INVX1_3/gnd DFFSR_23/S FILL
XFILL_1_DFFPOSX1_34 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_36_DFFSR_224 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_26_5_2 INVX1_3/gnd DFFSR_23/S FILL
XFILL_1_AND2X2_34 AND2X2_38/B DFFSR_59/S FILL
XFILL_12_DFFSR_123 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_6_BUFX2_30 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_26_DFFSR_227 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_2_AOI21X1_2 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_8_4_1 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_16_DFFSR_230 INVX1_67/gnd DFFSR_201/S FILL
XFILL_6_NAND3X1_149 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_6_6_2 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_43_DFFSR_52 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_8_DFFSR_117 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_32_DFFSR_92 BUFX2_99/A DFFSR_92/S FILL
XFILL_4_INVX1_86 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_49_DFFSR_148 INVX1_67/gnd DFFSR_175/S FILL
XNAND3X1_185 INVX1_157/Y OAI21X1_59/C OAI21X1_52/Y BUFX2_7/gnd NAND3X1_192/B DFFSR_216/S
+ NAND3X1
XFILL_39_DFFSR_151 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_16_DFFSR_42 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_2_DFFSR_227 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_3_BUFX2_77 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_29_DFFSR_154 BUFX2_99/A DFFSR_7/S FILL
XFILL_43_DFFSR_258 DFFSR_5/gnd DFFSR_5/S FILL
XNAND3X1_4 NAND3X1_4/A NAND3X1_4/B AND2X2_6/Y BUFX2_79/A NOR2X1_8/A DFFSR_7/S NAND3X1
XFILL_19_DFFSR_157 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_20_DFFPOSX1_42 INVX1_39/gnd DFFSR_34/S FILL
XFILL_33_DFFSR_261 BUFX2_77/gnd DFFSR_98/S FILL
XNOR2X1_39 NOR2X1_39/A NOR2X1_39/B OR2X2_6/gnd NOR2X1_39/Y DFFSR_92/S NOR2X1
XFILL_4_NAND3X1_1 BUFX2_98/A DFFSR_6/S FILL
XFILL_23_DFFSR_264 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_4_NAND3X1_245 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_40_DFFSR_99 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_4_NOR2X1_36 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_13_DFFSR_267 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_1_AND2X2_8 BUFX2_99/A DFFSR_7/S FILL
XFILL_7_OAI21X1_101 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_7_DFFSR_56 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_24_DFFSR_49 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_11_CLKBUF1_12 AND2X2_38/B DFFSR_23/S FILL
XFILL_5_DFFSR_154 BUFX2_99/A DFFSR_7/S FILL
XFILL_13_DFFSR_89 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_36_0_2 BUFX2_99/A DFFSR_92/S FILL
XFILL_5_NAND3X1_179 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_46_DFFSR_185 INVX1_39/gnd DFFSR_54/S FILL
XFILL_10_CLKBUF1_15 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_9_DFFSR_261 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_36_DFFSR_188 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_26_DFFSR_191 INVX1_67/gnd DFFSR_175/S FILL
XFILL_9_CLKBUF1_18 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_7_DFFSR_3 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_16_DFFSR_194 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_8_CLKBUF1_21 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_6_NAND3X1_113 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_7_CLKBUF1_24 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_10_DFFPOSX1_17 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_43_DFFSR_16 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_32_DFFSR_56 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_21_DFFSR_96 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_4_INVX1_50 BUFX2_98/A DFFSR_6/S FILL
XFILL_1_NOR2X1_73 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_6_CLKBUF1_27 INVX1_1/gnd DFFSR_97/S FILL
XFILL_49_DFFSR_112 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_5_CLKBUF1_30 BUFX2_77/gnd DFFSR_5/S FILL
XNAND3X1_149 INVX1_143/Y AOI22X1_20/A AOI21X1_15/B DFFSR_1/gnd AOI21X1_9/A DFFSR_1/S
+ NAND3X1
XFILL_39_DFFSR_115 INVX1_1/gnd DFFSR_97/S FILL
XCLKBUF1_27 BUFX2_6/Y INVX1_1/gnd CLKBUF1_27/Y DFFSR_97/S CLKBUF1
XFILL_2_DFFSR_191 INVX1_67/gnd DFFSR_175/S FILL
XFILL_4_CLKBUF1_33 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_5_OR2X2_3 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_3_BUFX2_41 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_29_DFFSR_118 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_43_DFFSR_222 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_3_CLKBUF1_36 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_8_AND2X2_32 AND2X2_38/B DFFSR_23/S FILL
XFILL_19_DFFSR_121 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_33_DFFSR_225 INVX1_67/gnd DFFSR_175/S FILL
XFILL_2_CLKBUF1_39 INVX1_1/gnd DFFSR_53/S FILL
XFILL_31_DFFSR_7 BUFX2_79/A DFFSR_7/S FILL
XFILL_23_DFFSR_228 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_1_CLKBUF1_42 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_4_NAND3X1_209 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_40_DFFSR_63 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_1_INVX1_97 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_0_DFFPOSX1_28 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_0_CLKBUF1_45 BUFX2_79/A DFFSR_7/S FILL
XFILL_13_DFFSR_231 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_7_DFFSR_20 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_24_DFFSR_13 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_5_DFFSR_118 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_13_DFFSR_53 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_0_BUFX2_88 INVX1_3/gnd DFFSR_23/S FILL
XFILL_46_DFFSR_149 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_5_NAND3X1_143 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_9_DFFSR_225 INVX1_67/gnd DFFSR_175/S FILL
XFILL_36_DFFSR_152 INVX1_1/gnd DFFSR_53/S FILL
XFILL_50_DFFSR_256 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_6_NOR2X1_1 BUFX2_99/A DFFSR_92/S FILL
XFILL_26_DFFSR_155 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_2_INVX1_202 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_40_DFFSR_259 BUFX2_79/A DFFSR_6/S FILL
XFILL_48_DFFSR_70 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_16_DFFSR_158 INVX1_3/gnd DFFSR_23/S FILL
XFILL_30_DFFSR_262 BUFX2_98/A DFFSR_32/S FILL
XFILL_1_NAND3X1_2 BUFX2_99/A DFFSR_7/S FILL
XFILL_20_DFFSR_265 INVX1_67/gnd DFFSR_175/S FILL
XFILL_19_DFFPOSX1_36 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_21_DFFSR_60 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_32_DFFSR_20 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_4_DFFSR_67 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_1_NOR2X1_37 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_27_6_0 INVX1_3/gnd DFFSR_79/S FILL
XFILL_10_DFFSR_268 OR2X2_1/gnd DFFSR_51/S FILL
XNAND3X1_113 DFFSR_191/D BUFX2_28/Y BUFX2_24/Y DFFSR_62/gnd NAND3X1_113/Y DFFSR_208/S
+ NAND3X1
XFILL_3_NAND3X1_239 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_2_DFFSR_155 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_43_DFFSR_186 BUFX2_99/A DFFSR_92/S FILL
XFILL_6_DFFSR_262 BUFX2_98/A DFFSR_32/S FILL
XFILL_33_DFFSR_189 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_23_DFFSR_192 INVX1_1/gnd DFFSR_97/S FILL
XFILL_4_NAND3X1_173 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_40_DFFSR_27 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_1_INVX1_61 INVX1_39/gnd DFFSR_54/S FILL
XFILL_29_DFFSR_67 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_13_DFFSR_195 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_9_DFFPOSX1_47 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_13_DFFSR_17 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_0_BUFX2_52 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_46_DFFSR_113 BUFX2_99/A DFFSR_92/S FILL
XFILL_5_NAND3X1_107 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_9_DFFSR_189 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_36_DFFSR_116 INVX1_3/gnd DFFSR_23/S FILL
XFILL_50_DFFSR_220 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_18_DFFSR_1 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_26_DFFSR_119 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_2_INVX1_166 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_40_DFFSR_223 INVX1_39/gnd DFFSR_34/S FILL
XFILL_37_DFFSR_74 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_5_AND2X2_33 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_48_DFFSR_34 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_16_DFFSR_122 BUFX2_79/A DFFSR_7/S FILL
XFILL_30_DFFSR_226 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_37_1_0 BUFX2_99/A DFFSR_7/S FILL
XFILL_6_AOI21X1_1 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_20_DFFSR_229 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_10_DFFSR_64 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_21_DFFSR_24 BUFX2_98/A DFFSR_6/S FILL
XFILL_4_DFFSR_31 BUFX2_79/A DFFSR_6/S FILL
XFILL_2_BUFX2_2 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_35_3_1 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_10_DFFSR_232 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_3_NAND3X1_203 INVX1_1/gnd DFFSR_97/S FILL
XFILL_9_OAI22X1_9 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_2_DFFSR_119 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_33_5_2 INVX1_1/gnd DFFSR_53/S FILL
XFILL_43_DFFSR_150 AND2X2_38/B DFFSR_23/S FILL
XFILL_45_DFFSR_81 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_6_DFFSR_226 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_33_DFFSR_153 INVX1_67/gnd DFFSR_201/S FILL
XFILL_47_DFFSR_257 INVX1_39/gnd DFFSR_34/S FILL
XFILL_23_DFFSR_156 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_4_NAND3X1_137 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_1_INVX1_25 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_1_DFFSR_78 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_37_DFFSR_260 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_29_DFFSR_31 BUFX2_79/A DFFSR_6/S FILL
XFILL_18_DFFSR_71 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_13_DFFSR_159 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_27_DFFSR_263 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_9_DFFPOSX1_11 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_6_NAND2X1_173 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_17_DFFSR_266 INVX1_67/gnd DFFSR_201/S FILL
XFILL_22_DFFPOSX1_3 INVX1_39/gnd DFFSR_34/S FILL
XFILL_0_BUFX2_16 BUFX2_98/A DFFSR_32/S FILL
XFILL_5_XOR2X1_8 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_21_DFFPOSX1_6 AND2X2_38/B DFFSR_23/S FILL
XFILL_9_DFFSR_153 INVX1_67/gnd DFFSR_201/S FILL
XFILL_20_DFFPOSX1_9 INVX1_67/gnd DFFSR_201/S FILL
XFILL_18_DFFPOSX1_30 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_50_DFFSR_184 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_2_INVX1_130 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_40_DFFSR_187 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_9_DFFSR_85 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_26_DFFSR_78 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_37_DFFSR_38 BUFX2_98/A DFFSR_6/S FILL
XFILL_2_NAND3X1_233 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_3_DFFSR_263 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_30_DFFSR_190 INVX1_39/gnd DFFSR_34/S FILL
XFILL_20_DFFSR_193 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_10_DFFSR_28 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_10_DFFSR_196 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_43_0_2 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_5_NOR2X1_72 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_3_NAND3X1_167 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_8_DFFPOSX1_41 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_43_DFFSR_114 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_45_DFFSR_45 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_34_DFFSR_85 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_6_DFFSR_190 INVX1_39/gnd DFFSR_34/S FILL
XFILL_33_DFFSR_117 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_47_DFFSR_221 AND2X2_38/B DFFSR_59/S FILL
XFILL_23_DFFSR_120 INVX1_3/gnd DFFSR_23/S FILL
XFILL_4_NAND3X1_101 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_37_DFFSR_224 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_1_DFFSR_42 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_18_DFFSR_35 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_2_AND2X2_34 AND2X2_38/B DFFSR_59/S FILL
XFILL_13_DFFSR_123 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_5_BUFX2_70 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_27_DFFSR_227 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_6_NAND2X1_137 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_3_AOI21X1_2 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_17_DFFSR_230 INVX1_67/gnd DFFSR_201/S FILL
XFILL_11_XOR2X1_5 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_9_DFFSR_117 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_42_DFFSR_92 BUFX2_99/A DFFSR_92/S FILL
XFILL_9_AOI21X1_62 INVX1_3/gnd DFFSR_23/S FILL
XNAND2X1_173 XOR2X1_9/A XOR2X1_9/B NOR3X1_6/gnd NAND2X1_173/Y DFFSR_79/S NAND2X1
XFILL_50_DFFSR_148 INVX1_67/gnd DFFSR_175/S FILL
XFILL_4_OAI21X1_119 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_27_DFFPOSX1_49 BUFX2_99/A DFFSR_92/S FILL
XFILL_8_AOI21X1_65 INVX1_3/gnd DFFSR_23/S FILL
XFILL_3_AND2X2_1 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_40_DFFSR_151 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_26_DFFSR_42 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_9_DFFSR_49 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_7_AOI21X1_68 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_15_DFFSR_82 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_2_NAND3X1_197 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_3_DFFSR_227 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_30_DFFSR_154 BUFX2_99/A DFFSR_7/S FILL
XFILL_6_AOI21X1_71 BUFX2_99/A DFFSR_92/S FILL
XFILL_44_DFFSR_258 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_20_DFFSR_157 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_34_DFFSR_261 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_5_NAND3X1_1 BUFX2_98/A DFFSR_6/S FILL
XAOI21X1_71 AOI21X1_71/A AOI21X1_71/B XNOR2X1_4/Y BUFX2_99/A NOR2X1_83/A DFFSR_92/S
+ AOI21X1
XFILL_10_DFFSR_160 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_24_DFFSR_264 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_50_DFFSR_99 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_3_NAND3X1_131 AND2X2_38/B DFFSR_59/S FILL
XFILL_5_NOR2X1_36 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_30_DFFSR_4 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_14_DFFSR_267 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_6_DFFSR_96 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_5_NAND2X1_167 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_6_DFFSR_154 BUFX2_99/A DFFSR_7/S FILL
XFILL_34_DFFSR_49 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_23_DFFSR_89 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_47_DFFSR_185 INVX1_39/gnd DFFSR_54/S FILL
XFILL_37_DFFSR_188 DFFSR_46/gnd DFFSR_54/S FILL
XBUFX2_74 BUFX2_74/A BUFX2_72/gnd dout[3] DFFSR_276/S BUFX2
XFILL_0_DFFSR_264 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_10_DFFPOSX1_3 INVX1_39/gnd DFFSR_34/S FILL
XFILL_5_BUFX2_34 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_27_DFFSR_191 INVX1_67/gnd DFFSR_175/S FILL
XFILL_34_6_0 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_17_DFFPOSX1_24 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_6_NAND2X1_101 INVX1_39/gnd DFFSR_54/S FILL
XFILL_17_DFFSR_194 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_1_NAND3X1_227 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_9_DFFPOSX1_6 AND2X2_38/B DFFSR_23/S FILL
XFILL_8_DFFPOSX1_9 INVX1_67/gnd DFFSR_201/S FILL
XFILL_42_DFFSR_56 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_31_DFFSR_96 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_3_INVX1_90 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_2_NOR2X1_73 OR2X2_3/gnd DFFSR_60/S FILL
XNAND2X1_137 DFFSR_62/S INVX1_195/A DFFSR_62/gnd OAI21X1_106/C DFFSR_62/S NAND2X1
XFILL_50_DFFSR_112 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_27_DFFPOSX1_13 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_8_AOI21X1_29 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_40_DFFSR_115 INVX1_1/gnd DFFSR_97/S FILL
XFILL_9_DFFSR_13 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_7_AOI21X1_32 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_2_NAND3X1_161 AND2X2_38/B DFFSR_23/S FILL
XFILL_15_DFFSR_46 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_3_DFFSR_191 INVX1_67/gnd DFFSR_175/S FILL
XFILL_30_DFFSR_118 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_2_BUFX2_81 BUFX2_79/A DFFSR_7/S FILL
XFILL_6_AOI21X1_35 INVX1_39/gnd DFFSR_54/S FILL
XFILL_44_DFFSR_222 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_20_DFFSR_121 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_7_DFFPOSX1_35 INVX1_39/gnd DFFSR_54/S FILL
XFILL_34_DFFSR_225 INVX1_67/gnd DFFSR_175/S FILL
XFILL_5_AOI21X1_38 DFFSR_28/gnd DFFSR_8/S FILL
XAOI21X1_35 OAI21X1_55/Y NAND2X1_91/Y INVX1_163/Y INVX1_39/gnd AOI21X1_35/Y DFFSR_54/S
+ AOI21X1
XFILL_10_DFFSR_124 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_4_AOI21X1_41 INVX1_39/gnd DFFSR_34/S FILL
XFILL_24_DFFSR_228 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_50_DFFSR_63 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_0_AOI21X1_3 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_3_AOI21X1_44 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_14_DFFSR_231 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_2_AOI21X1_47 INVX1_67/gnd DFFSR_175/S FILL
XFILL_6_DFFSR_60 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_5_NAND2X1_131 INVX1_3/gnd DFFSR_79/S FILL
XFILL_12_DFFSR_93 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_6_DFFSR_118 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_34_DFFSR_13 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_23_DFFSR_53 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_1_AOI21X1_50 INVX1_67/gnd DFFSR_175/S FILL
XFILL_47_DFFSR_149 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_44_1_0 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_0_AOI21X1_53 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_37_DFFSR_152 INVX1_1/gnd DFFSR_53/S FILL
XBUFX2_38 rst DFFSR_1/gnd BUFX2_38/Y DFFSR_1/S BUFX2
XFILL_0_DFFSR_228 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_27_DFFSR_155 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_3_OAI21X1_113 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_26_DFFPOSX1_43 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_41_DFFSR_259 BUFX2_79/A DFFSR_6/S FILL
XFILL_3_INVX1_202 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_42_3_1 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_17_DFFSR_158 INVX1_3/gnd DFFSR_23/S FILL
XFILL_8_OAI21X1_77 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_31_DFFSR_262 BUFX2_98/A DFFSR_32/S FILL
XFILL_1_NAND3X1_191 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_2_NAND3X1_2 BUFX2_99/A DFFSR_7/S FILL
XFILL_7_OAI21X1_80 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_6_NAND2X1_98 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_21_DFFSR_265 INVX1_67/gnd DFFSR_175/S FILL
XFILL_31_DFFSR_60 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_3_INVX1_54 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_42_DFFSR_20 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_40_5_2 BUFX2_98/A DFFSR_6/S FILL
XFILL_2_NOR2X1_37 BUFX2_7/gnd DFFSR_216/S FILL
XNAND2X1_101 NAND3X1_217/B NAND2X1_99/A INVX1_39/gnd INVX1_170/A DFFSR_54/S NAND2X1
XFILL_6_OAI21X1_83 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_11_DFFSR_268 OR2X2_1/gnd DFFSR_51/S FILL
XNAND2X1_98 NOR2X1_69/Y OAI21X1_63/Y OR2X2_6/gnd NAND2X1_98/Y DFFSR_53/S NAND2X1
XFILL_5_OAI21X1_86 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_15_DFFSR_10 DFFSR_5/gnd DFFSR_5/S FILL
XOAI21X1_83 AOI21X1_42/Y AOI21X1_35/Y AOI21X1_34/A DFFSR_34/gnd OAI21X1_83/Y DFFSR_1/S
+ OAI21X1
XFILL_2_NAND3X1_125 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_4_OAI21X1_89 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_3_DFFSR_155 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_2_BUFX2_45 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_44_DFFSR_186 BUFX2_99/A DFFSR_92/S FILL
XFILL_3_OAI21X1_92 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_7_DFFSR_262 BUFX2_98/A DFFSR_32/S FILL
XFILL_4_NAND2X1_161 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_34_DFFSR_189 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_2_OAI21X1_95 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_24_DFFSR_192 INVX1_1/gnd DFFSR_97/S FILL
XFILL_50_DFFSR_27 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_1_OAI21X1_98 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_39_DFFSR_67 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_14_DFFSR_195 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_3_1 INVX1_67/gnd DFFSR_201/S FILL
XFILL_2_AOI21X1_11 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_16_DFFPOSX1_18 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_6_DFFSR_24 BUFX2_98/A DFFSR_6/S FILL
XFILL_23_DFFSR_17 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_12_DFFSR_57 BUFX2_79/A DFFSR_6/S FILL
XFILL_1_AOI21X1_14 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_47_DFFSR_113 BUFX2_99/A DFFSR_92/S FILL
XFILL_0_NAND3X1_221 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_0_AOI21X1_17 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_37_DFFSR_116 INVX1_3/gnd DFFSR_23/S FILL
XFILL_51_DFFSR_220 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_5_NOR2X1_5 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_0_DFFSR_192 INVX1_1/gnd DFFSR_97/S FILL
XFILL_27_DFFSR_119 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_42_DFFSR_7 BUFX2_79/A DFFSR_7/S FILL
XFILL_9_OAI21X1_38 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_41_DFFSR_223 INVX1_39/gnd DFFSR_34/S FILL
XFILL_47_DFFSR_74 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_3_INVX1_166 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_6_AND2X2_33 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_50_0_2 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_17_DFFSR_122 BUFX2_79/A DFFSR_7/S FILL
XFILL_31_DFFSR_226 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_8_OAI21X1_41 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_1_NAND3X1_155 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_7_AOI21X1_1 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_6_NAND2X1_62 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_7_OAI21X1_44 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_21_DFFSR_229 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_31_DFFSR_24 BUFX2_98/A DFFSR_6/S FILL
XFILL_3_DFFSR_71 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_3_INVX1_18 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_6_DFFPOSX1_29 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_20_DFFSR_64 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_5_NAND2X1_65 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_6_OAI21X1_47 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_11_DFFSR_232 DFFSR_46/gnd DFFSR_54/S FILL
XNAND2X1_62 INVX1_133/A INVX1_175/A BUFX2_8/gnd INVX1_138/A DFFSR_81/S NAND2X1
XFILL_5_OAI21X1_50 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_4_NAND2X1_68 AND2X2_38/B DFFSR_23/S FILL
XOAI21X1_47 INVX1_145/Y INVX1_159/Y NAND2X1_71/Y DFFSR_34/gnd OAI21X1_47/Y DFFSR_1/S
+ OAI21X1
XFILL_3_DFFSR_119 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_3_NAND2X1_71 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_4_OAI21X1_53 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_7_XOR2X1_1 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_44_DFFSR_150 AND2X2_38/B DFFSR_23/S FILL
XFILL_15_DFFPOSX1_48 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_2_NAND2X1_74 AND2X2_38/B DFFSR_59/S FILL
XFILL_3_OAI21X1_56 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_7_DFFSR_226 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_34_DFFSR_153 INVX1_67/gnd DFFSR_201/S FILL
XFILL_4_NAND2X1_125 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_1_NAND2X1_77 AND2X2_38/B DFFSR_23/S FILL
XFILL_11_AOI22X1_25 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_48_DFFSR_257 INVX1_39/gnd DFFSR_34/S FILL
XFILL_2_OAI21X1_59 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_24_DFFSR_156 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_38_DFFSR_260 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_1_OAI21X1_62 INVX1_3/gnd DFFSR_79/S FILL
XFILL_0_NAND2X1_80 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_0_INVX1_203 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_0_INVX1_65 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_39_DFFSR_31 BUFX2_79/A DFFSR_6/S FILL
XFILL_10_AOI22X1_28 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_28_DFFSR_71 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_14_DFFSR_159 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_0_OAI21X1_65 INVX1_1/gnd DFFSR_53/S FILL
XFILL_16_1_1 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_28_DFFSR_263 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_2_OAI21X1_107 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_25_DFFPOSX1_37 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_18_DFFSR_266 INVX1_67/gnd DFFSR_201/S FILL
XFILL_12_DFFSR_21 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_14_3_2 INVX1_39/gnd DFFSR_54/S FILL
XFILL_0_NAND3X1_185 BUFX2_7/gnd DFFSR_216/S FILL
XNOR2X1_9 NOR2X1_9/A NOR2X1_9/B DFFSR_4/gnd NOR2X1_9/Y DFFSR_4/S NOR2X1
XFILL_3_NOR3X1_2 INVX1_1/gnd DFFSR_53/S FILL
XDFFSR_1 DFFSR_1/Q DFFSR_1/CLK DFFSR_1/R DFFSR_1/S DFFSR_1/D DFFSR_1/gnd DFFSR_1/S
+ DFFSR
XDFFSR_266 DFFSR_266/Q CLKBUF1_47/Y DFFSR_266/R DFFSR_201/S DFFSR_266/D INVX1_67/gnd
+ DFFSR_201/S DFFSR
XFILL_0_DFFSR_156 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_3_INVX1_130 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_41_DFFSR_187 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_36_DFFSR_78 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_47_DFFSR_38 BUFX2_98/A DFFSR_6/S FILL
XFILL_4_DFFSR_263 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_31_DFFSR_190 INVX1_39/gnd DFFSR_34/S FILL
XFILL_1_NAND3X1_119 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_6_NAND2X1_26 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_21_DFFSR_193 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_3_DFFSR_35 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_20_DFFSR_28 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_5_NAND2X1_29 INVX1_3/gnd DFFSR_23/S FILL
XFILL_6_OAI21X1_11 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_11_DFFSR_196 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_3_NAND2X1_155 BUFX2_79/A DFFSR_7/S FILL
XNAND2X1_26 DFFSR_40/Q AND2X2_5/Y DFFSR_8/gnd NAND2X1_26/Y DFFSR_8/S NAND2X1
XFILL_4_NAND2X1_32 INVX1_3/gnd DFFSR_79/S FILL
XFILL_5_OAI21X1_14 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_6_NOR2X1_72 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_8_6 BUFX2_7/gnd DFFSR_151/S FILL
XOAI21X1_11 INVX1_82/Y OAI21X1_9/B NAND2X1_41/Y XOR2X1_1/gnd NOR2X1_42/B DFFSR_208/S
+ OAI21X1
XFILL_3_NAND2X1_35 INVX1_67/gnd DFFSR_201/S FILL
XFILL_4_OAI21X1_17 DFFSR_46/gnd DFFSR_62/S FILL
XDFFPOSX1_29 DFFPOSX1_29/Q CLKBUF1_44/Y AOI21X1_57/Y BUFX2_72/gnd DFFSR_276/S DFFPOSX1
XFILL_44_DFFSR_114 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_41_6_0 BUFX2_98/A DFFSR_32/S FILL
XFILL_15_DFFPOSX1_12 AND2X2_38/B DFFSR_23/S FILL
XFILL_3_OAI21X1_20 AND2X2_38/B DFFSR_23/S FILL
XFILL_2_NAND2X1_38 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_29_DFFSR_1 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_44_DFFSR_85 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_7_DFFSR_190 INVX1_39/gnd DFFSR_34/S FILL
XFILL_34_DFFSR_117 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_2_OAI21X1_23 INVX1_67/gnd DFFSR_201/S FILL
XFILL_1_NAND2X1_41 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_48_DFFSR_221 AND2X2_38/B DFFSR_59/S FILL
XFILL_24_DFFSR_120 INVX1_3/gnd DFFSR_23/S FILL
XFILL_8_NAND3X1_97 AND2X2_38/B DFFSR_59/S FILL
XFILL_1_OAI21X1_26 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_38_DFFSR_224 BUFX2_7/gnd DFFSR_151/S FILL
XAOI21X1_5 OR2X2_1/B OR2X2_1/A NOR3X1_1/A INVX1_3/gnd NOR2X1_64/A DFFSR_23/S AOI21X1
XFILL_0_NAND2X1_44 INVX1_39/gnd DFFSR_34/S FILL
XFILL_28_DFFSR_35 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_0_INVX1_29 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_0_DFFSR_82 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_0_INVX1_167 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_17_DFFSR_75 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_3_AND2X2_34 AND2X2_38/B DFFSR_59/S FILL
XFILL_14_DFFSR_123 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_0_OAI21X1_29 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_28_DFFSR_227 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_4_AOI21X1_2 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_18_DFFSR_230 INVX1_67/gnd DFFSR_201/S FILL
XFILL_0_NAND3X1_149 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_9_NAND3X1_204 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_5_DFFPOSX1_23 NOR3X1_6/gnd DFFSR_91/S FILL
XDFFSR_230 DFFSR_238/D CLKBUF1_25/Y BUFX2_60/Y DFFSR_201/S DFFSR_222/Q INVX1_67/gnd
+ DFFSR_201/S DFFSR
XFILL_0_DFFSR_120 INVX1_3/gnd DFFSR_23/S FILL
XFILL_41_DFFSR_151 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_30_7 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_36_DFFSR_42 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_8_DFFSR_89 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_47_2 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_25_DFFSR_82 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_4_DFFSR_227 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_31_DFFSR_154 BUFX2_99/A DFFSR_7/S FILL
XFILL_45_DFFSR_258 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_4_AOI22X1_10 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_21_DFFSR_157 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_35_DFFSR_261 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_14_DFFPOSX1_42 INVX1_39/gnd DFFSR_34/S FILL
XFILL_3_AOI22X1_13 AND2X2_38/B DFFSR_23/S FILL
XFILL_6_NAND3X1_1 BUFX2_98/A DFFSR_6/S FILL
XFILL_3_NAND2X1_119 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_11_DFFSR_160 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_25_DFFSR_264 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_2_AOI22X1_16 BUFX2_77/gnd DFFSR_5/S FILL
XINVX1_3 INVX1_3/A INVX1_3/gnd INVX1_3/Y DFFSR_79/S INVX1
XFILL_6_NOR2X1_36 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_51_1_0 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_15_DFFSR_267 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_17_NOR3X1_6 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_1_AOI22X1_19 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_0_AOI22X1_22 INVX1_3/gnd DFFSR_79/S FILL
XFILL_10_OAI22X1_40 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_44_DFFSR_49 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_33_DFFSR_89 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_1_OAI21X1_101 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_7_DFFSR_154 BUFX2_99/A DFFSR_7/S FILL
XFILL_24_DFFPOSX1_31 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_49_3_1 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_48_DFFSR_185 INVX1_39/gnd DFFSR_54/S FILL
XFILL_8_NAND3X1_61 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_9_OAI22X1_43 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_38_DFFSR_188 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_0_INVX1_131 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_8_NAND3X1_234 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_17_DFFSR_39 INVX1_3/gnd DFFSR_79/S FILL
XFILL_0_DFFSR_46 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_4_BUFX2_74 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_47_5_2 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_1_DFFSR_264 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_7_NAND3X1_64 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_8_OAI22X1_46 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_28_DFFSR_191 INVX1_67/gnd DFFSR_175/S FILL
XFILL_6_NAND3X1_67 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_7_OAI22X1_49 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_18_DFFSR_194 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_5_NAND3X1_70 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_6_OAI22X1_52 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_0_NAND3X1_113 DFFSR_62/gnd DFFSR_208/S FILL
XNAND3X1_67 BUFX2_90/A AND2X2_16/Y BUFX2_34/Y XOR2X1_1/gnd AND2X2_19/A DFFSR_151/S
+ NAND3X1
XFILL_10_XOR2X1_9 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_4_NAND3X1_73 INVX1_1/gnd DFFSR_97/S FILL
XFILL_41_DFFSR_96 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_3_NOR2X1_73 OR2X2_3/gnd DFFSR_60/S FILL
XOAI22X1_52 AOI21X1_44/Y AOI21X1_45/Y OAI21X1_84/Y AND2X2_40/Y DFFSR_28/gnd OAI22X1_52/Y
+ DFFSR_3/S OAI22X1
XFILL_3_NAND3X1_76 INVX1_1/gnd DFFSR_53/S FILL
XFILL_2_NAND2X1_149 OR2X2_2/gnd DFFSR_216/S FILL
XDFFSR_194 DFFSR_194/Q CLKBUF1_6/Y BUFX2_70/Y DFFSR_81/S DFFSR_194/D DFFSR_1/gnd DFFSR_81/S
+ DFFSR
XFILL_2_AND2X2_5 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_41_DFFSR_115 INVX1_1/gnd DFFSR_97/S FILL
XFILL_2_NAND3X1_79 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_8_DFFSR_53 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_14_DFFSR_86 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_25_DFFSR_46 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_4_DFFSR_191 INVX1_67/gnd DFFSR_175/S FILL
XFILL_31_DFFSR_118 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_15_4_0 INVX1_39/gnd DFFSR_34/S FILL
XFILL_1_NAND3X1_82 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_45_DFFSR_222 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_21_DFFSR_121 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_0_NAND3X1_85 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_35_DFFSR_225 INVX1_67/gnd DFFSR_175/S FILL
XFILL_0_AND2X2_35 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_11_DFFSR_124 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_13_6_1 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_25_DFFSR_228 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_1_AOI21X1_3 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_20_DFFSR_8 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_15_DFFSR_231 DFFSR_46/gnd DFFSR_62/S FILL
XINVX1_87 INVX1_87/A OR2X2_2/gnd INVX1_87/Y DFFSR_175/S INVX1
XFILL_22_DFFSR_93 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_44_DFFSR_13 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_33_DFFSR_53 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_7_DFFSR_118 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_48_DFFSR_149 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_8_NAND3X1_25 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_4_BUFX2_9 AND2X2_38/B DFFSR_59/S FILL
XFILL_38_DFFSR_152 INVX1_1/gnd DFFSR_53/S FILL
XFILL_8_NAND3X1_198 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_0_DFFSR_10 DFFSR_5/gnd DFFSR_5/S FILL
XINVX1_205 BUFX2_77/A BUFX2_99/A INVX1_205/Y DFFSR_92/S INVX1
XFILL_7_NAND3X1_28 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_8_OAI22X1_10 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_4_BUFX2_38 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_1_DFFSR_228 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_28_DFFSR_155 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_4_DFFPOSX1_17 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_42_DFFSR_259 BUFX2_79/A DFFSR_6/S FILL
XFILL_1_NAND2X1_179 INVX1_1/gnd DFFSR_97/S FILL
XFILL_4_INVX1_202 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_6_NAND3X1_31 BUFX2_79/A DFFSR_6/S FILL
XFILL_7_OAI22X1_13 INVX1_1/gnd DFFSR_53/S FILL
XFILL_18_DFFSR_158 INVX1_3/gnd DFFSR_23/S FILL
XFILL_5_NAND3X1_34 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_32_DFFSR_262 BUFX2_98/A DFFSR_32/S FILL
XFILL_41_DFFSR_4 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_3_NAND3X1_2 BUFX2_99/A DFFSR_7/S FILL
XFILL_6_OAI22X1_16 AND2X2_38/B DFFSR_59/S FILL
XNAND3X1_31 NAND3X1_31/A NAND3X1_31/B AOI22X1_4/Y BUFX2_79/A NOR2X1_17/B DFFSR_6/S
+ NAND3X1
XFILL_22_DFFSR_265 INVX1_67/gnd DFFSR_175/S FILL
XFILL_2_INVX1_94 INVX1_67/gnd DFFSR_201/S FILL
XFILL_5_OAI22X1_19 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_4_NAND3X1_37 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_41_DFFSR_60 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_3_NOR2X1_37 BUFX2_7/gnd DFFSR_216/S FILL
XOAI22X1_16 INVX1_38/Y OAI22X1_7/B INVX1_39/Y OAI22X1_7/D AND2X2_38/B NOR2X1_21/B
+ DFFSR_59/S OAI22X1
XFILL_13_DFFPOSX1_36 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_12_DFFSR_268 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_4_OAI22X1_22 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_3_NAND3X1_40 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_2_NAND2X1_113 OR2X2_4/gnd DFFSR_3/S FILL
XDFFSR_158 INVX1_102/A CLKBUF1_22/Y BUFX2_61/Y DFFSR_23/S DFFSR_158/D INVX1_3/gnd
+ DFFSR_23/S DFFSR
XFILL_2_NAND3X1_43 BUFX2_99/A DFFSR_7/S FILL
XFILL_3_OAI22X1_25 INVX1_39/gnd DFFSR_54/S FILL
XFILL_8_DFFSR_17 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_25_DFFSR_10 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_14_DFFSR_50 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_4_DFFSR_155 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_1_BUFX2_85 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_1_NAND3X1_46 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_2_OAI22X1_28 INVX1_3/gnd DFFSR_23/S FILL
XFILL_45_DFFSR_186 BUFX2_99/A DFFSR_92/S FILL
XFILL_23_1_1 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_0_NAND3X1_49 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_8_DFFSR_262 BUFX2_98/A DFFSR_32/S FILL
XFILL_1_OAI22X1_31 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_35_DFFSR_189 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_5_0_0 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_23_DFFPOSX1_25 BUFX2_79/A DFFSR_6/S FILL
XFILL_0_OAI22X1_34 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_25_DFFSR_192 INVX1_1/gnd DFFSR_97/S FILL
XFILL_21_3_2 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_49_DFFSR_67 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_7_NAND3X1_228 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_15_DFFSR_195 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_3_2_1 INVX1_67/gnd DFFSR_175/S FILL
XFILL_3_DFFPOSX1_47 XOR2X1_4/gnd DFFSR_91/S FILL
XINVX1_51 INVX1_51/A DFFSR_28/gnd INVX1_51/Y DFFSR_8/S INVX1
XFILL_33_DFFSR_17 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_5_DFFSR_64 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_22_DFFSR_57 BUFX2_79/A DFFSR_6/S FILL
XFILL_11_DFFSR_97 INVX1_1/gnd DFFSR_97/S FILL
XFILL_0_NOR2X1_74 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_1_4_2 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_48_DFFSR_113 BUFX2_99/A DFFSR_92/S FILL
XFILL_38_DFFSR_116 INVX1_3/gnd DFFSR_23/S FILL
XFILL_8_NAND3X1_162 BUFX2_8/gnd DFFSR_51/S FILL
XINVX1_169 INVX1_169/A INVX1_39/gnd INVX1_169/Y DFFSR_34/S INVX1
XFILL_1_DFFSR_192 INVX1_1/gnd DFFSR_97/S FILL
XFILL_28_DFFSR_119 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_1_NAND2X1_143 INVX1_67/gnd DFFSR_201/S FILL
XFILL_42_DFFSR_223 INVX1_39/gnd DFFSR_34/S FILL
XFILL_4_INVX1_166 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_7_AND2X2_33 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_18_DFFSR_122 BUFX2_79/A DFFSR_7/S FILL
XFILL_32_DFFSR_226 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_8_AOI21X1_1 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_22_DFFSR_229 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_41_DFFSR_24 BUFX2_98/A DFFSR_6/S FILL
XFILL_2_INVX1_58 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_30_DFFSR_64 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_48_6_0 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_12_DFFSR_232 DFFSR_46/gnd DFFSR_54/S FILL
XDFFSR_122 BUFX2_83/A CLKBUF1_40/Y BUFX2_49/Y DFFSR_7/S INVX1_16/A BUFX2_79/A DFFSR_7/S
+ DFFSR
XFILL_14_DFFSR_14 INVX1_1/gnd DFFSR_53/S FILL
XFILL_4_DFFSR_119 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_1_NAND3X1_10 BUFX2_79/A DFFSR_6/S FILL
XFILL_1_BUFX2_49 INVX1_1/gnd DFFSR_97/S FILL
XFILL_45_DFFSR_150 AND2X2_38/B DFFSR_23/S FILL
XFILL_0_NAND3X1_13 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_8_DFFSR_226 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_35_DFFSR_153 INVX1_67/gnd DFFSR_201/S FILL
XFILL_8_DFFSR_7 BUFX2_79/A DFFSR_7/S FILL
XFILL_49_DFFSR_257 INVX1_39/gnd DFFSR_34/S FILL
XFILL_9_OAI21X1_114 AND2X2_38/B DFFSR_59/S FILL
XFILL_25_DFFSR_156 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_39_DFFSR_260 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_1_INVX1_203 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_49_DFFSR_31 BUFX2_79/A DFFSR_6/S FILL
XFILL_38_DFFSR_71 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_7_NAND3X1_192 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_15_DFFSR_159 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_29_DFFSR_263 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_0_NAND3X1_3 BUFX2_99/A DFFSR_92/S FILL
XFILL_3_DFFPOSX1_11 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_19_DFFSR_266 INVX1_67/gnd DFFSR_201/S FILL
XINVX1_15 DFFSR_18/D BUFX2_98/A INVX1_15/Y DFFSR_32/S INVX1
XDFFSR_68 DFFSR_76/D DFFSR_7/CLK DFFSR_9/R DFFSR_6/S DFFSR_68/D BUFX2_98/A DFFSR_6/S
+ DFFSR
XFILL_0_NAND2X1_173 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_5_DFFSR_28 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_22_DFFSR_21 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_11_DFFSR_61 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_0_NOR2X1_38 INVX1_3/gnd DFFSR_79/S FILL
XFILL_8_NAND3X1_126 DFFSR_62/gnd DFFSR_62/S FILL
XINVX1_133 INVX1_133/A OR2X2_1/gnd INVX1_133/Y DFFSR_51/S INVX1
XFILL_4_NOR2X1_9 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_1_DFFSR_156 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_12_DFFPOSX1_30 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_1_NAND2X1_107 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_42_DFFSR_187 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_4_INVX1_130 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_46_DFFSR_78 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_5_DFFSR_263 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_32_DFFSR_190 INVX1_39/gnd DFFSR_34/S FILL
XFILL_22_DFFSR_193 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_2_INVX1_22 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_2_DFFSR_75 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_30_DFFSR_28 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_19_DFFSR_68 BUFX2_98/A DFFSR_6/S FILL
XFILL_12_DFFSR_196 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_22_DFFPOSX1_19 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_1_BUFX2_13 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_6_NAND3X1_222 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_54_5_2 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_6_XOR2X1_5 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_45_DFFSR_114 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_2_DFFPOSX1_41 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_8_DFFSR_190 INVX1_39/gnd DFFSR_34/S FILL
XFILL_35_DFFSR_117 BUFX2_77/gnd DFFSR_98/S FILL
XAND2X2_37 BUFX2_59/Y AND2X2_37/B XOR2X1_4/gnd AND2X2_37/Y DFFSR_97/S AND2X2
XFILL_49_DFFSR_221 AND2X2_38/B DFFSR_59/S FILL
XFILL_25_DFFSR_120 INVX1_3/gnd DFFSR_23/S FILL
XFILL_39_DFFSR_224 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_38_DFFSR_35 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_1_INVX1_167 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_27_DFFSR_75 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_4_AND2X2_34 AND2X2_38/B DFFSR_59/S FILL
XFILL_15_DFFSR_123 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_7_NAND3X1_156 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_29_DFFSR_227 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_5_AOI21X1_2 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_19_DFFSR_230 INVX1_67/gnd DFFSR_201/S FILL
XDFFSR_32 DFFSR_24/D DFFSR_8/CLK DFFSR_2/R DFFSR_32/S DFFSR_8/Q OR2X2_4/gnd DFFSR_32/S
+ DFFSR
XFILL_0_NAND2X1_137 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_11_DFFSR_25 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_22_4_0 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_2_NOR3X1_6 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_1_DFFSR_120 INVX1_3/gnd DFFSR_23/S FILL
XFILL_42_DFFSR_151 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_21_DFFPOSX1_49 BUFX2_99/A DFFSR_92/S FILL
XFILL_20_6_1 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_35_DFFSR_82 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_46_DFFSR_42 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_5_DFFSR_227 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_32_DFFSR_154 BUFX2_99/A DFFSR_7/S FILL
XFILL_2_5_0 INVX1_67/gnd DFFSR_201/S FILL
XFILL_46_DFFSR_258 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_22_DFFSR_157 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_2_DFFSR_39 INVX1_3/gnd DFFSR_79/S FILL
XFILL_36_DFFSR_261 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_19_DFFSR_32 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_7_NAND3X1_1 BUFX2_98/A DFFSR_6/S FILL
XFILL_6_BUFX2_67 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_12_DFFSR_160 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_26_DFFSR_264 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_8_OAI21X1_108 INVX1_1/gnd DFFSR_53/S FILL
XFILL_16_DFFSR_267 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_6_NAND3X1_186 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_20_CLKBUF1_22 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_12_XOR2X1_2 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_19_DFFSR_5 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_19_CLKBUF1_25 INVX1_67/gnd DFFSR_201/S FILL
XFILL_43_DFFSR_89 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_8_DFFSR_154 BUFX2_99/A DFFSR_7/S FILL
XFILL_18_CLKBUF1_28 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_49_DFFSR_185 INVX1_39/gnd DFFSR_54/S FILL
XNAND3X1_222 NAND2X1_90/A NAND3X1_217/B NAND3X1_216/Y DFFSR_46/gnd AOI21X1_40/A DFFSR_54/S
+ NAND3X1
XFILL_17_CLKBUF1_31 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_39_DFFSR_188 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_1_INVX1_131 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_27_DFFSR_39 INVX1_3/gnd DFFSR_79/S FILL
XFILL_16_DFFSR_79 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_2_DFFSR_264 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_7_NAND3X1_120 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_16_CLKBUF1_34 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_29_DFFSR_191 INVX1_67/gnd DFFSR_175/S FILL
XFILL_3_BUFX2_6 BUFX2_79/A DFFSR_6/S FILL
XFILL_11_DFFPOSX1_24 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_15_CLKBUF1_37 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_19_DFFSR_194 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_0_NAND2X1_101 INVX1_39/gnd DFFSR_54/S FILL
XNOR2X1_76 NOR2X1_76/A NOR2X1_76/B INVX1_3/gnd NOR2X1_76/Y DFFSR_79/S NOR2X1
XFILL_14_CLKBUF1_40 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_4_NOR2X1_73 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_30_1_1 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_13_CLKBUF1_43 AND2X2_38/B DFFSR_23/S FILL
XFILL_40_DFFSR_1 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_12_CLKBUF1_46 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_42_DFFSR_115 INVX1_1/gnd DFFSR_97/S FILL
XFILL_21_DFFPOSX1_13 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_7_DFFSR_93 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_24_DFFSR_86 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_11_CLKBUF1_49 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_35_DFFSR_46 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_5_DFFSR_191 INVX1_67/gnd DFFSR_175/S FILL
XFILL_28_3_2 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_32_DFFSR_118 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_46_DFFSR_222 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_5_NAND3X1_216 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_22_DFFSR_121 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_36_DFFSR_225 INVX1_67/gnd DFFSR_175/S FILL
XFILL_1_DFFPOSX1_35 INVX1_39/gnd DFFSR_54/S FILL
XFILL_1_AND2X2_35 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_12_DFFSR_124 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_6_BUFX2_31 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_26_DFFSR_228 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_2_AOI21X1_3 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_8_4_2 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_16_DFFSR_231 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_6_NAND3X1_150 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_43_DFFSR_53 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_32_DFFSR_93 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_8_DFFSR_118 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_49_DFFSR_149 BUFX2_72/gnd DFFSR_276/S FILL
XNAND3X1_186 INVX1_157/A OAI21X1_53/Y OAI21X1_54/Y BUFX2_7/gnd NAND3X1_192/C DFFSR_151/S
+ NAND3X1
XFILL_39_DFFSR_152 INVX1_1/gnd DFFSR_53/S FILL
XFILL_16_DFFSR_43 BUFX2_98/A DFFSR_6/S FILL
XFILL_2_DFFSR_228 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_3_BUFX2_78 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_29_DFFSR_155 OR2X2_1/gnd DFFSR_59/S FILL
XNAND3X1_5 DFFSR_9/Q BUFX2_22/Y BUFX2_11/Y BUFX2_99/A NAND3X1_7/A DFFSR_7/S NAND3X1
XFILL_43_DFFSR_259 BUFX2_79/A DFFSR_6/S FILL
XFILL_20_DFFPOSX1_43 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_19_DFFSR_158 INVX1_3/gnd DFFSR_23/S FILL
XFILL_33_DFFSR_262 BUFX2_98/A DFFSR_32/S FILL
XFILL_4_NAND3X1_2 BUFX2_99/A DFFSR_7/S FILL
XNOR2X1_40 NOR2X1_40/A NOR2X1_40/B NOR3X1_6/gnd NOR2X1_40/Y DFFSR_91/S NOR2X1
XFILL_23_DFFSR_265 INVX1_67/gnd DFFSR_175/S FILL
XFILL_4_NAND3X1_246 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_51_DFFSR_60 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_4_NOR2X1_37 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_13_DFFSR_268 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_12_CLKBUF1_10 INVX1_67/gnd DFFSR_201/S FILL
XFILL_7_OAI21X1_102 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_1_AND2X2_9 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_11_CLKBUF1_13 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_35_DFFSR_10 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_24_DFFSR_50 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_13_DFFSR_90 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_7_DFFSR_57 BUFX2_79/A DFFSR_6/S FILL
XFILL_5_DFFSR_155 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_10_CLKBUF1_16 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_46_DFFSR_186 BUFX2_99/A DFFSR_92/S FILL
XFILL_5_NAND3X1_180 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_9_DFFSR_262 BUFX2_98/A DFFSR_32/S FILL
XFILL_36_DFFSR_189 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_26_DFFSR_192 INVX1_1/gnd DFFSR_97/S FILL
XFILL_9_CLKBUF1_19 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_7_DFFSR_4 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_8_CLKBUF1_22 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_16_DFFSR_195 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_6_NAND3X1_114 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_7_CLKBUF1_25 INVX1_67/gnd DFFSR_201/S FILL
XFILL_10_DFFPOSX1_18 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_43_DFFSR_17 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_32_DFFSR_57 BUFX2_79/A DFFSR_6/S FILL
XFILL_21_DFFSR_97 INVX1_1/gnd DFFSR_97/S FILL
XFILL_6_CLKBUF1_28 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_1_NOR2X1_74 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_49_DFFSR_113 BUFX2_99/A DFFSR_92/S FILL
XFILL_5_CLKBUF1_31 BUFX2_72/gnd DFFSR_201/S FILL
XNAND3X1_150 AOI21X1_12/B AOI21X1_12/A AOI21X1_8/Y DFFSR_1/gnd NAND3X1_152/C DFFSR_1/S
+ NAND3X1
XFILL_39_DFFSR_116 INVX1_3/gnd DFFSR_23/S FILL
XCLKBUF1_28 BUFX2_1/Y OR2X2_4/gnd DFFSR_2/CLK DFFSR_3/S CLKBUF1
XFILL_4_CLKBUF1_34 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_5_OR2X2_4 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_2_DFFSR_192 INVX1_1/gnd DFFSR_97/S FILL
XFILL_3_BUFX2_42 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_29_DFFSR_119 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_43_DFFSR_223 INVX1_39/gnd DFFSR_34/S FILL
XFILL_3_CLKBUF1_37 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_8_AND2X2_33 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_19_DFFSR_122 BUFX2_79/A DFFSR_7/S FILL
XFILL_33_DFFSR_226 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_2_CLKBUF1_40 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_31_DFFSR_8 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_9_AOI21X1_1 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_1_CLKBUF1_43 AND2X2_38/B DFFSR_23/S FILL
XFILL_23_DFFSR_229 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_4_NAND3X1_210 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_40_DFFSR_64 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_51_DFFSR_24 BUFX2_98/A DFFSR_6/S FILL
XFILL_1_INVX1_98 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_0_DFFPOSX1_29 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_13_DFFSR_232 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_0_CLKBUF1_46 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_16_1 INVX1_39/gnd DFFSR_34/S FILL
XFILL_7_DFFSR_21 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_24_DFFSR_14 INVX1_1/gnd DFFSR_53/S FILL
XFILL_13_DFFSR_54 INVX1_39/gnd DFFSR_54/S FILL
XFILL_5_DFFSR_119 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_0_BUFX2_89 INVX1_1/gnd DFFSR_97/S FILL
XFILL_46_DFFSR_150 AND2X2_38/B DFFSR_23/S FILL
XFILL_5_NAND3X1_144 AND2X2_38/B DFFSR_59/S FILL
XFILL_9_DFFSR_226 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_36_DFFSR_153 INVX1_67/gnd DFFSR_201/S FILL
XFILL_6_NOR2X1_2 INVX1_1/gnd DFFSR_97/S FILL
XFILL_50_DFFSR_257 INVX1_39/gnd DFFSR_34/S FILL
XFILL_26_DFFSR_156 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_2_INVX1_203 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_40_DFFSR_260 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_48_DFFSR_71 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_29_4_0 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_16_DFFSR_159 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_30_DFFSR_263 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_1_NAND3X1_3 BUFX2_99/A DFFSR_92/S FILL
XFILL_20_DFFSR_266 INVX1_67/gnd DFFSR_201/S FILL
XFILL_32_DFFSR_21 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_4_INVX1_15 BUFX2_98/A DFFSR_32/S FILL
XFILL_4_DFFSR_68 BUFX2_98/A DFFSR_6/S FILL
XFILL_19_DFFPOSX1_37 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_21_DFFSR_61 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_27_6_1 INVX1_3/gnd DFFSR_79/S FILL
XFILL_1_NOR2X1_38 INVX1_3/gnd DFFSR_79/S FILL
XFILL_10_DFFSR_269 INVX1_67/gnd DFFSR_201/S FILL
XFILL_9_5_0 XOR2X1_1/gnd DFFSR_208/S FILL
XNAND3X1_114 DFFSR_135/Q AND2X2_18/B BUFX2_28/Y XOR2X1_1/gnd AND2X2_25/B DFFSR_208/S
+ NAND3X1
XFILL_3_NAND3X1_240 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_2_DFFSR_156 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_43_DFFSR_187 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_6_DFFSR_263 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_33_DFFSR_190 INVX1_39/gnd DFFSR_34/S FILL
XFILL_23_DFFSR_193 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_4_NAND3X1_174 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_40_DFFSR_28 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_29_DFFSR_68 BUFX2_98/A DFFSR_6/S FILL
XFILL_1_INVX1_62 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_13_DFFSR_196 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_0_CLKBUF1_10 INVX1_67/gnd DFFSR_201/S FILL
XFILL_9_DFFPOSX1_48 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_13_DFFSR_18 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_0_BUFX2_53 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_46_DFFSR_114 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_5_NAND3X1_108 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_9_DFFSR_190 INVX1_39/gnd DFFSR_34/S FILL
XFILL_36_DFFSR_117 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_50_DFFSR_221 AND2X2_38/B DFFSR_59/S FILL
XFILL_18_DFFSR_2 BUFX2_79/A DFFSR_7/S FILL
XFILL_26_DFFSR_120 INVX1_3/gnd DFFSR_23/S FILL
XFILL_40_DFFSR_224 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_48_DFFSR_35 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_2_INVX1_167 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_5_AND2X2_34 AND2X2_38/B DFFSR_59/S FILL
XFILL_37_DFFSR_75 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_16_DFFSR_123 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_30_DFFSR_227 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_37_1_1 BUFX2_99/A DFFSR_7/S FILL
XFILL_6_AOI21X1_2 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_20_DFFSR_230 INVX1_67/gnd DFFSR_201/S FILL
XFILL_4_DFFSR_32 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_21_DFFSR_25 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_10_DFFSR_65 BUFX2_79/A DFFSR_7/S FILL
XFILL_2_BUFX2_3 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_10_DFFSR_233 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_35_3_2 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_3_NAND3X1_204 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_2_DFFSR_120 INVX1_3/gnd DFFSR_23/S FILL
XFILL_43_DFFSR_151 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_45_DFFSR_82 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_6_DFFSR_227 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_33_DFFSR_154 BUFX2_99/A DFFSR_7/S FILL
XFILL_47_DFFSR_258 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_4_NAND3X1_138 INVX1_67/gnd DFFSR_201/S FILL
XFILL_23_DFFSR_157 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_18_DFFSR_72 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_37_DFFSR_261 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_29_DFFSR_32 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_1_INVX1_26 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_1_DFFSR_79 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_8_NAND3X1_1 BUFX2_98/A DFFSR_6/S FILL
XFILL_13_DFFSR_160 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_27_DFFSR_264 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_9_DFFPOSX1_12 AND2X2_38/B DFFSR_23/S FILL
XFILL_23_DFFPOSX1_1 INVX1_39/gnd DFFSR_34/S FILL
XFILL_6_NAND2X1_174 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_17_DFFSR_267 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_22_DFFPOSX1_4 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_0_BUFX2_17 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_5_XOR2X1_9 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_21_DFFPOSX1_7 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_9_DFFSR_154 BUFX2_99/A DFFSR_7/S FILL
XFILL_18_DFFPOSX1_31 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_50_DFFSR_185 INVX1_39/gnd DFFSR_54/S FILL
XFILL_2_INVX1_131 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_9_DFFSR_86 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_40_DFFSR_188 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_26_DFFSR_79 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_37_DFFSR_39 INVX1_3/gnd DFFSR_79/S FILL
XFILL_3_DFFSR_264 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_2_NAND3X1_234 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_30_DFFSR_191 INVX1_67/gnd DFFSR_175/S FILL
XFILL_20_DFFSR_194 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_10_DFFSR_29 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_10_DFFSR_197 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_5_NOR2X1_73 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_3_NAND3X1_168 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_43_DFFSR_115 INVX1_1/gnd DFFSR_97/S FILL
XFILL_8_DFFPOSX1_42 INVX1_39/gnd DFFSR_34/S FILL
XFILL_34_DFFSR_86 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_45_DFFSR_46 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_6_DFFSR_191 INVX1_67/gnd DFFSR_175/S FILL
XFILL_33_DFFSR_118 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_47_DFFSR_222 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_23_DFFSR_121 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_4_NAND3X1_102 INVX1_3/gnd DFFSR_23/S FILL
XFILL_37_DFFSR_225 INVX1_67/gnd DFFSR_175/S FILL
XFILL_18_DFFSR_36 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_1_DFFSR_43 BUFX2_98/A DFFSR_6/S FILL
XFILL_2_AND2X2_35 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_13_DFFSR_124 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_5_BUFX2_71 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_27_DFFSR_228 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_6_NAND2X1_138 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_3_AOI21X1_3 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_17_DFFSR_231 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_6_DFFSR_1 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_11_XOR2X1_6 BUFX2_99/A DFFSR_7/S FILL
XFILL_42_DFFSR_93 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_9_DFFSR_118 OR2X2_3/gnd DFFSR_60/S FILL
XNAND2X1_174 NOR2X1_80/A NOR2X1_80/B XOR2X1_4/gnd AOI21X1_66/B DFFSR_91/S NAND2X1
XFILL_50_DFFSR_149 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_8_AOI21X1_66 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_27_DFFPOSX1_50 INVX1_1/gnd DFFSR_53/S FILL
XFILL_3_AND2X2_2 BUFX2_99/A DFFSR_7/S FILL
XFILL_40_DFFSR_152 INVX1_1/gnd DFFSR_53/S FILL
XFILL_9_DFFSR_50 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_26_DFFSR_43 BUFX2_98/A DFFSR_6/S FILL
XFILL_7_AOI21X1_69 INVX1_1/gnd DFFSR_97/S FILL
XFILL_15_DFFSR_83 INVX1_3/gnd DFFSR_79/S FILL
XFILL_2_NAND3X1_198 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_3_DFFSR_228 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_30_DFFSR_155 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_44_DFFSR_259 BUFX2_79/A DFFSR_6/S FILL
XFILL_20_DFFSR_158 INVX1_3/gnd DFFSR_23/S FILL
XFILL_4_OR2X2_1 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_34_DFFSR_262 BUFX2_98/A DFFSR_32/S FILL
XFILL_5_NAND3X1_2 BUFX2_99/A DFFSR_7/S FILL
XFILL_10_DFFSR_161 INVX1_67/gnd DFFSR_175/S FILL
XFILL_24_DFFSR_265 INVX1_67/gnd DFFSR_175/S FILL
XFILL_5_NOR2X1_37 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_3_NAND3X1_132 AND2X2_38/B DFFSR_23/S FILL
XFILL_30_DFFSR_5 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_14_DFFSR_268 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_45_DFFSR_10 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_34_DFFSR_50 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_5_NAND2X1_168 BUFX2_79/A DFFSR_6/S FILL
XFILL_6_DFFSR_97 INVX1_1/gnd DFFSR_97/S FILL
XFILL_23_DFFSR_90 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_6_DFFSR_155 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_36_4_0 BUFX2_99/A DFFSR_92/S FILL
XFILL_47_DFFSR_186 BUFX2_99/A DFFSR_92/S FILL
XFILL_11_DFFPOSX1_1 INVX1_39/gnd DFFSR_34/S FILL
XFILL_37_DFFSR_189 BUFX2_8/gnd DFFSR_51/S FILL
XBUFX2_75 BUFX2_75/A BUFX2_72/gnd dout[4] DFFSR_276/S BUFX2
XFILL_0_DFFSR_265 INVX1_67/gnd DFFSR_175/S FILL
XFILL_17_DFFPOSX1_25 BUFX2_79/A DFFSR_6/S FILL
XFILL_34_6_1 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_5_BUFX2_35 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_10_DFFPOSX1_4 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_27_DFFSR_192 INVX1_1/gnd DFFSR_97/S FILL
XFILL_6_NAND2X1_102 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_17_DFFSR_195 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_1_NAND3X1_228 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_9_DFFPOSX1_7 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_42_DFFSR_57 BUFX2_79/A DFFSR_6/S FILL
XFILL_31_DFFSR_97 INVX1_1/gnd DFFSR_97/S FILL
XFILL_3_INVX1_91 AND2X2_38/B DFFSR_23/S FILL
XNAND2X1_138 DFFSR_7/S INVX1_196/A OR2X2_6/gnd OAI21X1_107/C DFFSR_92/S NAND2X1
XFILL_2_NOR2X1_74 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_50_DFFSR_113 BUFX2_99/A DFFSR_92/S FILL
XFILL_8_AOI21X1_30 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_27_DFFPOSX1_14 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_40_DFFSR_116 INVX1_3/gnd DFFSR_23/S FILL
XFILL_9_DFFSR_14 INVX1_1/gnd DFFSR_53/S FILL
XFILL_15_DFFSR_47 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_7_AOI21X1_33 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_3_DFFSR_192 INVX1_1/gnd DFFSR_97/S FILL
XFILL_2_NAND3X1_162 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_2_BUFX2_82 INVX1_1/gnd DFFSR_97/S FILL
XFILL_30_DFFSR_119 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_6_AOI21X1_36 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_44_DFFSR_223 INVX1_39/gnd DFFSR_34/S FILL
XFILL_9_AND2X2_33 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_7_DFFPOSX1_36 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_20_DFFSR_122 BUFX2_79/A DFFSR_7/S FILL
XFILL_5_AOI21X1_39 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_34_DFFSR_226 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_10_DFFSR_125 DFFSR_5/gnd DFFSR_5/S FILL
XAOI21X1_36 AOI21X1_36/A AOI21X1_36/B INVX1_173/Y BUFX2_77/gnd OAI21X1_80/A DFFSR_98/S
+ AOI21X1
XFILL_4_AOI21X1_42 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_24_DFFSR_229 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_50_DFFSR_64 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_0_AOI21X1_4 BUFX2_98/A DFFSR_32/S FILL
XFILL_3_AOI21X1_45 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_14_DFFSR_232 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_2_AOI21X1_48 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_5_NAND2X1_132 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_6_DFFSR_61 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_34_DFFSR_14 INVX1_1/gnd DFFSR_53/S FILL
XFILL_6_DFFSR_119 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_12_DFFSR_94 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_1_AOI21X1_51 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_23_DFFSR_54 INVX1_39/gnd DFFSR_54/S FILL
XFILL_47_DFFSR_150 AND2X2_38/B DFFSR_23/S FILL
XFILL_44_1_1 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_0_AOI21X1_54 AND2X2_38/B DFFSR_59/S FILL
XFILL_37_DFFSR_153 INVX1_67/gnd DFFSR_201/S FILL
XBUFX2_39 rst BUFX2_7/gnd BUFX2_39/Y DFFSR_151/S BUFX2
XFILL_0_DFFSR_229 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_27_DFFSR_156 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_3_OAI21X1_114 AND2X2_38/B DFFSR_59/S FILL
XFILL_3_INVX1_203 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_26_DFFPOSX1_44 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_41_DFFSR_260 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_42_3_2 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_17_DFFSR_159 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_1_NAND3X1_192 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_8_OAI21X1_78 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_31_DFFSR_263 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_2_NAND3X1_3 BUFX2_99/A DFFSR_92/S FILL
XFILL_21_DFFSR_266 INVX1_67/gnd DFFSR_201/S FILL
XFILL_7_OAI21X1_81 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_6_NAND2X1_99 INVX1_39/gnd DFFSR_54/S FILL
XFILL_31_DFFSR_61 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_3_INVX1_55 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_42_DFFSR_21 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_2_NOR2X1_38 INVX1_3/gnd DFFSR_79/S FILL
XNAND2X1_102 XNOR2X1_1/B XNOR2X1_1/A OR2X2_1/gnd INVX1_172/A DFFSR_51/S NAND2X1
XFILL_6_OAI21X1_84 BUFX2_98/A DFFSR_6/S FILL
XFILL_11_DFFSR_269 INVX1_67/gnd DFFSR_201/S FILL
XNAND2X1_99 NAND2X1_99/A NAND2X1_99/B INVX1_39/gnd NAND2X1_99/Y DFFSR_54/S NAND2X1
XFILL_5_OAI21X1_87 BUFX2_79/A DFFSR_7/S FILL
XOAI21X1_84 INVX1_180/Y AND2X2_40/A INVX1_131/Y BUFX2_98/A OAI21X1_84/Y DFFSR_6/S
+ OAI21X1
XFILL_15_DFFSR_11 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_3_DFFSR_156 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_2_NAND3X1_126 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_4_OAI21X1_90 BUFX2_98/A DFFSR_32/S FILL
XFILL_2_BUFX2_46 BUFX2_98/A DFFSR_6/S FILL
XFILL_44_DFFSR_187 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_3_OAI21X1_93 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_10_2_0 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_7_DFFSR_263 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_4_NAND2X1_162 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_34_DFFSR_190 INVX1_39/gnd DFFSR_34/S FILL
XFILL_2_OAI21X1_96 AND2X2_38/B DFFSR_59/S FILL
XFILL_24_DFFSR_193 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_1_OAI21X1_99 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_50_DFFSR_28 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_39_DFFSR_68 BUFX2_98/A DFFSR_6/S FILL
XFILL_14_DFFSR_196 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_3_2 INVX1_67/gnd DFFSR_201/S FILL
XFILL_2_AOI21X1_12 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_16_DFFPOSX1_19 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_6_DFFSR_25 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_23_DFFSR_18 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_12_DFFSR_58 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_1_AOI21X1_15 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_47_DFFSR_114 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_0_NAND3X1_222 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_0_AOI21X1_18 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_37_DFFSR_117 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_0_DFFSR_193 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_5_NOR2X1_6 BUFX2_98/A DFFSR_6/S FILL
XFILL_27_DFFSR_120 INVX1_3/gnd DFFSR_23/S FILL
XFILL_42_DFFSR_8 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_41_DFFSR_224 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_3_INVX1_167 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_6_AND2X2_34 AND2X2_38/B DFFSR_59/S FILL
XFILL_47_DFFSR_75 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_17_DFFSR_123 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_8_OAI21X1_42 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_31_DFFSR_227 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_1_NAND3X1_156 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_7_AOI21X1_2 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_21_DFFSR_230 INVX1_67/gnd DFFSR_201/S FILL
XFILL_6_NAND2X1_63 AND2X2_38/B DFFSR_59/S FILL
XFILL_7_OAI21X1_45 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_3_DFFSR_72 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_31_DFFSR_25 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_20_DFFSR_65 BUFX2_79/A DFFSR_7/S FILL
XFILL_3_INVX1_19 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_6_DFFPOSX1_30 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_6_OAI21X1_48 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_5_NAND2X1_66 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_11_DFFSR_233 OR2X2_2/gnd DFFSR_175/S FILL
XNAND2X1_63 BUFX2_57/Y INVX1_145/A AND2X2_38/B NOR2X1_65/B DFFSR_59/S NAND2X1
XFILL_4_NAND2X1_69 INVX1_3/gnd DFFSR_23/S FILL
XFILL_5_OAI21X1_51 DFFSR_62/gnd DFFSR_208/S FILL
XOAI21X1_48 INVX1_134/Y INVX1_150/Y AND2X2_36/Y BUFX2_8/gnd OAI21X1_48/Y DFFSR_81/S
+ OAI21X1
XFILL_3_DFFSR_120 INVX1_3/gnd DFFSR_23/S FILL
XFILL_3_NAND2X1_72 AND2X2_38/B DFFSR_59/S FILL
XFILL_2_BUFX2_10 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_4_OAI21X1_54 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_7_XOR2X1_2 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_44_DFFSR_151 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_15_DFFPOSX1_49 BUFX2_99/A DFFSR_92/S FILL
XFILL_2_NAND2X1_75 INVX1_3/gnd DFFSR_79/S FILL
XFILL_3_OAI21X1_57 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_7_DFFSR_227 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_4_NAND2X1_126 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_34_DFFSR_154 BUFX2_99/A DFFSR_7/S FILL
XFILL_1_NAND2X1_78 AND2X2_38/B DFFSR_23/S FILL
XFILL_2_OAI21X1_60 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_48_DFFSR_258 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_11_AOI22X1_26 INVX1_1/gnd DFFSR_97/S FILL
XFILL_24_DFFSR_157 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_1_OAI21X1_63 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_0_NAND2X1_81 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_0_INVX1_66 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_0_INVX1_204 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_38_DFFSR_261 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_39_DFFSR_32 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_10_AOI22X1_29 INVX1_1/gnd DFFSR_53/S FILL
XFILL_28_DFFSR_72 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_9_NAND3X1_1 BUFX2_98/A DFFSR_6/S FILL
XFILL_14_DFFSR_160 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_16_1_2 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_28_DFFSR_264 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_0_OAI21X1_66 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_2_OAI21X1_108 INVX1_1/gnd DFFSR_53/S FILL
XFILL_25_DFFPOSX1_38 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_18_DFFSR_267 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_12_DFFSR_22 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_0_NAND3X1_186 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_9_NAND3X1_241 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_3_NOR3X1_3 BUFX2_7/gnd DFFSR_216/S FILL
XDFFSR_2 DFFSR_2/Q DFFSR_2/CLK DFFSR_2/R DFFSR_7/S DFFSR_2/D BUFX2_79/A DFFSR_7/S
+ DFFSR
XFILL_51_DFFSR_185 INVX1_39/gnd DFFSR_54/S FILL
XFILL_0_DFFSR_157 XOR2X1_1/gnd DFFSR_151/S FILL
XDFFSR_267 INVX1_192/A CLKBUF1_44/Y DFFSR_266/R DFFSR_208/S DFFSR_267/D XOR2X1_1/gnd
+ DFFSR_208/S DFFSR
XFILL_3_INVX1_131 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_41_DFFSR_188 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_36_DFFSR_79 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_47_DFFSR_39 INVX1_3/gnd DFFSR_79/S FILL
XFILL_4_DFFSR_264 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_31_DFFSR_191 INVX1_67/gnd DFFSR_175/S FILL
XFILL_1_NAND3X1_120 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_6_NAND2X1_27 AND2X2_38/B DFFSR_23/S FILL
XFILL_21_DFFSR_194 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_20_DFFSR_29 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_3_DFFSR_36 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_5_NAND2X1_30 AND2X2_38/B DFFSR_23/S FILL
XFILL_3_NAND2X1_156 AND2X2_38/B DFFSR_59/S FILL
XFILL_6_OAI21X1_12 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_11_DFFSR_197 XOR2X1_4/gnd DFFSR_97/S FILL
XNAND2X1_27 BUFX2_25/Y AND2X2_15/Y AND2X2_38/B OAI22X1_43/D DFFSR_23/S NAND2X1
XFILL_43_4_0 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_4_NAND2X1_33 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_5_OAI21X1_15 INVX1_3/gnd DFFSR_79/S FILL
XFILL_6_NOR2X1_73 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_8_7 BUFX2_7/gnd DFFSR_151/S FILL
XOAI21X1_12 INVX1_89/Y OAI21X1_9/B NAND2X1_43/Y OR2X2_1/gnd NOR2X1_45/B DFFSR_51/S
+ OAI21X1
XFILL_3_NAND2X1_36 INVX1_3/gnd DFFSR_79/S FILL
XFILL_4_OAI21X1_18 INVX1_39/gnd DFFSR_34/S FILL
XDFFPOSX1_30 NAND2X1_153/B CLKBUF1_46/Y AOI21X1_53/Y BUFX2_77/gnd DFFSR_98/S DFFPOSX1
XFILL_44_DFFSR_115 INVX1_1/gnd DFFSR_97/S FILL
XFILL_41_6_1 BUFX2_98/A DFFSR_32/S FILL
XFILL_29_DFFSR_2 BUFX2_79/A DFFSR_7/S FILL
XFILL_44_DFFSR_86 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_2_NAND2X1_39 BUFX2_98/A DFFSR_6/S FILL
XFILL_3_OAI21X1_21 AND2X2_38/B DFFSR_59/S FILL
XFILL_15_DFFPOSX1_13 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_7_DFFSR_191 INVX1_67/gnd DFFSR_175/S FILL
XFILL_34_DFFSR_118 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_2_OAI21X1_24 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_1_NAND2X1_42 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_48_DFFSR_222 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_24_DFFSR_121 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_8_NAND3X1_98 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_1_OAI21X1_27 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_0_NAND2X1_45 INVX1_39/gnd DFFSR_34/S FILL
XFILL_38_DFFSR_225 INVX1_67/gnd DFFSR_175/S FILL
XFILL_0_INVX1_168 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_0_INVX1_30 INVX1_1/gnd DFFSR_53/S FILL
XFILL_0_DFFSR_83 INVX1_3/gnd DFFSR_79/S FILL
XAOI21X1_6 AOI21X1_6/A AOI21X1_6/B BUFX2_38/Y DFFSR_1/gnd AOI21X1_6/Y DFFSR_81/S AOI21X1
XFILL_28_DFFSR_36 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_17_DFFSR_76 BUFX2_79/A DFFSR_7/S FILL
XFILL_3_AND2X2_35 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_14_DFFSR_124 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_0_OAI21X1_30 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_28_DFFSR_228 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_4_AOI21X1_3 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_18_DFFSR_231 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_0_NAND3X1_150 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_51_DFFSR_149 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_0_DFFSR_121 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_5_DFFPOSX1_24 BUFX2_8/gnd DFFSR_51/S FILL
XDFFSR_231 DFFSR_231/Q CLKBUF1_29/Y BUFX2_66/Y DFFSR_62/S DFFSR_231/D DFFSR_46/gnd
+ DFFSR_62/S DFFSR
XFILL_41_DFFSR_152 INVX1_1/gnd DFFSR_53/S FILL
XFILL_8_DFFSR_90 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_36_DFFSR_43 BUFX2_98/A DFFSR_6/S FILL
XFILL_25_DFFSR_83 INVX1_3/gnd DFFSR_79/S FILL
XFILL_47_3 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_4_DFFSR_228 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_31_DFFSR_155 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_45_DFFSR_259 BUFX2_79/A DFFSR_6/S FILL
XFILL_4_AOI22X1_11 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_21_DFFSR_158 INVX1_3/gnd DFFSR_23/S FILL
XFILL_14_DFFPOSX1_43 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_35_DFFSR_262 BUFX2_98/A DFFSR_32/S FILL
XFILL_3_AOI22X1_14 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_11_DFFSR_161 INVX1_67/gnd DFFSR_175/S FILL
XFILL_6_NAND3X1_2 BUFX2_99/A DFFSR_7/S FILL
XFILL_3_NAND2X1_120 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_25_DFFSR_265 INVX1_67/gnd DFFSR_175/S FILL
XFILL_2_AOI22X1_17 NOR3X1_6/gnd DFFSR_79/S FILL
XINVX1_4 OR2X2_1/A BUFX2_99/A INVX1_4/Y DFFSR_7/S INVX1
XFILL_6_NOR2X1_37 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_51_1_1 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_15_DFFSR_268 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_1_AOI22X1_20 INVX1_39/gnd DFFSR_34/S FILL
XFILL_0_AOI22X1_23 INVX1_39/gnd DFFSR_34/S FILL
XFILL_10_OAI22X1_41 INVX1_39/gnd DFFSR_54/S FILL
XFILL_44_DFFSR_50 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_1_OAI21X1_102 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_33_DFFSR_90 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_7_DFFSR_155 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_24_DFFPOSX1_32 INVX1_67/gnd DFFSR_201/S FILL
XFILL_49_3_2 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_48_DFFSR_186 BUFX2_99/A DFFSR_92/S FILL
XFILL_8_NAND3X1_62 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_9_OAI22X1_44 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_8_NAND3X1_235 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_0_DFFSR_47 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_0_INVX1_132 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_38_DFFSR_189 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_17_DFFSR_40 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_4_BUFX2_75 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_1_DFFSR_265 INVX1_67/gnd DFFSR_175/S FILL
XFILL_8_OAI22X1_47 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_7_NAND3X1_65 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_28_DFFSR_192 INVX1_1/gnd DFFSR_97/S FILL
XFILL_6_NAND3X1_68 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_7_OAI22X1_50 INVX1_3/gnd DFFSR_23/S FILL
XFILL_18_DFFSR_195 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_5_NAND3X1_71 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_0_NAND3X1_114 XOR2X1_1/gnd DFFSR_208/S FILL
XNAND3X1_68 NAND2X1_37/Y NAND3X1_68/B AND2X2_19/Y BUFX2_7/gnd NOR2X1_37/A DFFSR_216/S
+ NAND3X1
XFILL_4_NAND3X1_74 INVX1_1/gnd DFFSR_97/S FILL
XFILL_41_DFFSR_97 INVX1_1/gnd DFFSR_97/S FILL
XFILL_3_NOR2X1_74 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_17_2_0 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_3_NAND3X1_77 DFFSR_5/gnd DFFSR_5/S FILL
XDFFSR_195 DFFSR_195/Q CLKBUF1_11/Y BUFX2_69/Y DFFSR_62/S DFFSR_195/D DFFSR_46/gnd
+ DFFSR_62/S DFFSR
XFILL_2_NAND2X1_150 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_2_AND2X2_6 BUFX2_99/A DFFSR_7/S FILL
XFILL_2_NAND3X1_80 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_41_DFFSR_116 INVX1_3/gnd DFFSR_23/S FILL
XFILL_25_DFFSR_47 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_8_DFFSR_54 INVX1_39/gnd DFFSR_54/S FILL
XFILL_14_DFFSR_87 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_4_DFFSR_192 INVX1_1/gnd DFFSR_97/S FILL
XFILL_15_4_1 INVX1_39/gnd DFFSR_34/S FILL
XFILL_1_NAND3X1_83 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_31_DFFSR_119 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_45_DFFSR_223 INVX1_39/gnd DFFSR_34/S FILL
XFILL_21_DFFSR_122 BUFX2_79/A DFFSR_7/S FILL
XFILL_0_NAND3X1_86 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_35_DFFSR_226 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_0_AND2X2_36 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_11_DFFSR_125 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_13_6_2 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_25_DFFSR_229 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_1_AOI21X1_4 BUFX2_98/A DFFSR_32/S FILL
XFILL_20_DFFSR_9 BUFX2_79/A DFFSR_6/S FILL
XFILL_15_DFFSR_232 DFFSR_46/gnd DFFSR_54/S FILL
XINVX1_88 INVX1_88/A OR2X2_2/gnd INVX1_88/Y DFFSR_216/S INVX1
XFILL_44_DFFSR_14 INVX1_1/gnd DFFSR_53/S FILL
XFILL_7_DFFSR_119 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_22_DFFSR_94 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_33_DFFSR_54 INVX1_39/gnd DFFSR_54/S FILL
XFILL_48_DFFSR_150 AND2X2_38/B DFFSR_23/S FILL
XFILL_8_NAND3X1_26 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_38_DFFSR_153 INVX1_67/gnd DFFSR_201/S FILL
XINVX1_206 BUFX2_78/A INVX1_1/gnd INVX1_206/Y DFFSR_53/S INVX1
XFILL_8_NAND3X1_199 INVX1_1/gnd DFFSR_97/S FILL
XFILL_0_DFFSR_11 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_4_BUFX2_39 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_7_NAND3X1_29 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_8_OAI22X1_11 BUFX2_99/A DFFSR_92/S FILL
XFILL_1_DFFSR_229 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_28_DFFSR_156 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_4_DFFPOSX1_18 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_4_INVX1_203 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_42_DFFSR_260 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_1_NAND2X1_180 INVX1_1/gnd DFFSR_97/S FILL
XFILL_7_OAI22X1_14 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_6_NAND3X1_32 BUFX2_79/A DFFSR_7/S FILL
XFILL_18_DFFSR_159 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_32_DFFSR_263 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_5_NAND3X1_35 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_6_OAI22X1_17 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_41_DFFSR_5 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_3_NAND3X1_3 BUFX2_99/A DFFSR_92/S FILL
XNAND3X1_32 NOR2X1_15/Y NOR2X1_16/Y NOR2X1_17/Y BUFX2_79/A XOR2X1_11/A DFFSR_7/S NAND3X1
XFILL_22_DFFSR_266 INVX1_67/gnd DFFSR_201/S FILL
XFILL_5_OAI22X1_20 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_4_NAND3X1_38 BUFX2_98/A DFFSR_32/S FILL
XFILL_2_INVX1_95 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_41_DFFSR_61 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_3_NOR2X1_38 INVX1_3/gnd DFFSR_79/S FILL
XFILL_13_DFFPOSX1_37 BUFX2_72/gnd DFFSR_201/S FILL
XOAI22X1_17 INVX1_40/Y OAI22X1_2/B INVX1_41/Y OAI22X1_2/D DFFSR_4/gnd NOR2X1_21/A
+ DFFSR_98/S OAI22X1
XFILL_12_DFFSR_269 INVX1_67/gnd DFFSR_201/S FILL
XFILL_4_OAI22X1_23 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_3_NAND3X1_41 OR2X2_6/gnd DFFSR_92/S FILL
XDFFSR_159 DFFSR_151/D CLKBUF1_20/Y BUFX2_69/Y DFFSR_208/S DFFSR_135/Q DFFSR_62/gnd
+ DFFSR_208/S DFFSR
XFILL_2_NAND2X1_114 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_2_NAND3X1_44 BUFX2_99/A DFFSR_7/S FILL
XFILL_3_OAI22X1_26 INVX1_39/gnd DFFSR_54/S FILL
XFILL_8_DFFSR_18 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_25_DFFSR_11 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_4_DFFSR_156 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_14_DFFSR_51 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_1_NAND3X1_47 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_1_BUFX2_86 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_2_OAI22X1_29 INVX1_3/gnd DFFSR_79/S FILL
XFILL_23_1_2 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_45_DFFSR_187 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_0_NAND3X1_50 BUFX2_98/A DFFSR_6/S FILL
XFILL_8_DFFSR_263 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_1_OAI22X1_32 INVX1_39/gnd DFFSR_54/S FILL
XFILL_35_DFFSR_190 INVX1_39/gnd DFFSR_34/S FILL
XFILL_5_0_1 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_23_DFFPOSX1_26 AND2X2_38/B DFFSR_23/S FILL
XFILL_0_OAI22X1_35 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_25_DFFSR_193 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_49_DFFSR_68 BUFX2_98/A DFFSR_6/S FILL
XFILL_15_DFFSR_196 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_7_NAND3X1_229 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_3_2_2 INVX1_67/gnd DFFSR_175/S FILL
XFILL_3_DFFPOSX1_48 XOR2X1_4/gnd DFFSR_97/S FILL
XINVX1_52 DFFSR_16/D DFFSR_8/gnd INVX1_52/Y DFFSR_8/S INVX1
XFILL_5_DFFSR_65 BUFX2_79/A DFFSR_7/S FILL
XFILL_22_DFFSR_58 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_11_DFFSR_98 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_33_DFFSR_18 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_0_NOR2X1_75 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_48_DFFSR_114 NOR3X1_6/gnd DFFSR_91/S FILL
XINVX1_170 INVX1_170/A DFFSR_28/gnd INVX1_170/Y DFFSR_8/S INVX1
XFILL_38_DFFSR_117 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_8_NAND3X1_163 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_1_DFFSR_193 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_28_DFFSR_120 INVX1_3/gnd DFFSR_23/S FILL
XFILL_42_DFFSR_224 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_4_INVX1_167 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_1_NAND2X1_144 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_7_AND2X2_34 AND2X2_38/B DFFSR_59/S FILL
XFILL_50_4_0 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_18_DFFSR_123 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_32_DFFSR_227 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_8_AOI21X1_2 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_22_DFFSR_230 INVX1_67/gnd DFFSR_201/S FILL
XFILL_41_DFFSR_25 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_30_DFFSR_65 BUFX2_79/A DFFSR_7/S FILL
XFILL_2_INVX1_59 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_48_6_1 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_12_DFFSR_233 OR2X2_2/gnd DFFSR_175/S FILL
XDFFSR_123 BUFX2_84/A CLKBUF1_27/Y BUFX2_49/Y DFFSR_97/S INVX1_23/A XOR2X1_4/gnd DFFSR_97/S
+ DFFSR
XFILL_14_DFFSR_15 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_4_DFFSR_120 INVX1_3/gnd DFFSR_23/S FILL
XFILL_1_BUFX2_50 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_1_NAND3X1_11 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_45_DFFSR_151 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_8_DFFSR_227 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_0_NAND3X1_14 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_8_DFFSR_8 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_35_DFFSR_154 BUFX2_99/A DFFSR_7/S FILL
XFILL_49_DFFSR_258 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_25_DFFSR_157 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_1_INVX1_204 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_39_DFFSR_261 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_49_DFFSR_32 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_38_DFFSR_72 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_15_DFFSR_160 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_7_NAND3X1_193 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_29_DFFSR_264 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_0_NAND3X1_4 BUFX2_79/A DFFSR_7/S FILL
XFILL_3_DFFPOSX1_12 AND2X2_38/B DFFSR_23/S FILL
XFILL_0_NAND2X1_174 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_5_DFFSR_29 BUFX2_77/gnd DFFSR_5/S FILL
XDFFSR_69 DFFSR_69/Q DFFSR_57/CLK DFFSR_9/R DFFSR_32/S DFFSR_13/Q BUFX2_98/A DFFSR_32/S
+ DFFSR
XINVX1_16 INVX1_16/A BUFX2_99/A INVX1_16/Y DFFSR_7/S INVX1
XFILL_19_DFFSR_267 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_22_DFFSR_22 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_11_DFFSR_62 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_0_NOR2X1_39 OR2X2_6/gnd DFFSR_92/S FILL
XINVX1_134 AND2X2_35/A INVX1_3/gnd INVX1_134/Y DFFSR_79/S INVX1
XFILL_8_NAND3X1_127 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_1_DFFSR_157 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_12_DFFPOSX1_31 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_1_NAND2X1_108 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_42_DFFSR_188 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_46_DFFSR_79 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_5_DFFSR_264 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_32_DFFSR_191 INVX1_67/gnd DFFSR_175/S FILL
XFILL_22_DFFSR_194 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_30_DFFSR_29 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_2_DFFSR_76 BUFX2_79/A DFFSR_7/S FILL
XFILL_2_INVX1_23 BUFX2_99/A DFFSR_7/S FILL
XFILL_19_DFFSR_69 BUFX2_98/A DFFSR_32/S FILL
XFILL_12_DFFSR_197 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_22_DFFPOSX1_20 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_1_BUFX2_14 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_6_NAND3X1_223 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_6_XOR2X1_6 BUFX2_99/A DFFSR_7/S FILL
XFILL_45_DFFSR_115 INVX1_1/gnd DFFSR_97/S FILL
XFILL_8_DFFSR_191 INVX1_67/gnd DFFSR_175/S FILL
XFILL_2_DFFPOSX1_42 INVX1_39/gnd DFFSR_34/S FILL
XFILL_35_DFFSR_118 OR2X2_3/gnd DFFSR_60/S FILL
XAND2X2_38 INVX1_133/A AND2X2_38/B AND2X2_38/B XNOR2X1_1/B DFFSR_59/S AND2X2
XFILL_49_DFFSR_222 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_25_DFFSR_121 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_39_DFFSR_225 INVX1_67/gnd DFFSR_175/S FILL
XFILL_1_INVX1_168 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_38_DFFSR_36 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_27_DFFSR_76 BUFX2_79/A DFFSR_7/S FILL
XFILL_4_AND2X2_35 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_15_DFFSR_124 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_7_NAND3X1_157 INVX1_3/gnd DFFSR_23/S FILL
XFILL_29_DFFSR_228 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_24_2_0 AND2X2_38/B DFFSR_59/S FILL
XFILL_5_AOI21X1_3 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_0_NAND2X1_138 OR2X2_6/gnd DFFSR_92/S FILL
XDFFSR_33 DFFSR_41/D CLKBUF1_7/Y DFFSR_3/R DFFSR_32/S INVX1_7/A BUFX2_98/A DFFSR_32/S
+ DFFSR
XFILL_19_DFFSR_231 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_11_DFFSR_26 BUFX2_79/A DFFSR_6/S FILL
XFILL_22_4_1 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_4_3_0 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_1_DFFSR_121 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_21_DFFPOSX1_50 INVX1_1/gnd DFFSR_53/S FILL
XFILL_42_DFFSR_152 INVX1_1/gnd DFFSR_53/S FILL
XFILL_20_6_2 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_46_DFFSR_43 BUFX2_98/A DFFSR_6/S FILL
XFILL_35_DFFSR_83 INVX1_3/gnd DFFSR_79/S FILL
XFILL_5_DFFSR_228 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_32_DFFSR_155 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_2_5_1 INVX1_67/gnd DFFSR_201/S FILL
XFILL_46_DFFSR_259 BUFX2_79/A DFFSR_6/S FILL
XFILL_22_DFFSR_158 INVX1_3/gnd DFFSR_23/S FILL
XFILL_2_DFFSR_40 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_36_DFFSR_262 BUFX2_98/A DFFSR_32/S FILL
XFILL_19_DFFSR_33 BUFX2_98/A DFFSR_32/S FILL
XFILL_7_NAND3X1_2 BUFX2_99/A DFFSR_7/S FILL
XFILL_12_DFFSR_161 INVX1_67/gnd DFFSR_175/S FILL
XFILL_6_BUFX2_68 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_26_DFFSR_265 INVX1_67/gnd DFFSR_175/S FILL
XFILL_8_OAI21X1_109 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_21_CLKBUF1_20 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_16_DFFSR_268 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_6_NAND3X1_187 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_12_XOR2X1_3 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_19_DFFSR_6 BUFX2_79/A DFFSR_6/S FILL
XFILL_19_CLKBUF1_26 INVX1_1/gnd DFFSR_53/S FILL
XFILL_43_DFFSR_90 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_8_DFFSR_155 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_49_DFFSR_186 BUFX2_99/A DFFSR_92/S FILL
XFILL_18_CLKBUF1_29 XOR2X1_4/gnd DFFSR_91/S FILL
XNAND3X1_223 AOI21X1_25/Y NAND3X1_218/Y NAND3X1_219/Y DFFSR_46/gnd AOI21X1_40/B DFFSR_54/S
+ NAND3X1
XFILL_1_INVX1_132 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_39_DFFSR_189 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_17_CLKBUF1_32 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_27_DFFSR_40 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_16_DFFSR_80 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_2_DFFSR_265 INVX1_67/gnd DFFSR_175/S FILL
XFILL_7_NAND3X1_121 INVX1_1/gnd DFFSR_97/S FILL
XFILL_16_CLKBUF1_35 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_29_DFFSR_192 INVX1_1/gnd DFFSR_97/S FILL
XFILL_3_BUFX2_7 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_11_DFFPOSX1_25 BUFX2_79/A DFFSR_6/S FILL
XFILL_0_NAND2X1_102 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_15_CLKBUF1_38 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_19_DFFSR_195 DFFSR_46/gnd DFFSR_62/S FILL
XNOR2X1_77 NOR2X1_77/A NOR2X1_77/B INVX1_39/gnd NOR2X1_77/Y DFFSR_34/S NOR2X1
XFILL_14_CLKBUF1_41 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_30_1_2 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_13_CLKBUF1_44 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_4_NOR2X1_74 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_40_DFFSR_2 BUFX2_79/A DFFSR_7/S FILL
XFILL_12_CLKBUF1_47 BUFX2_98/A DFFSR_32/S FILL
XFILL_21_DFFPOSX1_14 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_42_DFFSR_116 INVX1_3/gnd DFFSR_23/S FILL
XFILL_35_DFFSR_47 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_7_DFFSR_94 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_24_DFFSR_87 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_5_DFFSR_192 INVX1_1/gnd DFFSR_97/S FILL
XFILL_32_DFFSR_119 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_46_DFFSR_223 INVX1_39/gnd DFFSR_34/S FILL
XFILL_5_NAND3X1_217 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_22_DFFSR_122 BUFX2_79/A DFFSR_7/S FILL
XFILL_1_DFFPOSX1_36 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_36_DFFSR_226 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_1_AND2X2_36 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_12_DFFSR_125 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_6_BUFX2_32 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_26_DFFSR_229 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_2_AOI21X1_4 BUFX2_98/A DFFSR_32/S FILL
XFILL_16_DFFSR_232 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_6_NAND3X1_151 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_4_INVX1_88 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_8_DFFSR_119 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_32_DFFSR_94 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_43_DFFSR_54 INVX1_39/gnd DFFSR_54/S FILL
XFILL_49_DFFSR_150 AND2X2_38/B DFFSR_23/S FILL
XNAND3X1_187 NOR3X1_5/B NAND3X1_192/B NAND3X1_192/C BUFX2_7/gnd NAND3X1_187/Y DFFSR_216/S
+ NAND3X1
XFILL_39_DFFSR_153 INVX1_67/gnd DFFSR_201/S FILL
XFILL_16_DFFSR_44 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_2_DFFSR_229 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_29_DFFSR_156 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_3_BUFX2_79 BUFX2_79/A DFFSR_7/S FILL
XFILL_43_DFFSR_260 BUFX2_77/gnd DFFSR_5/S FILL
XNAND3X1_6 DFFSR_73/D BUFX2_16/Y NOR2X1_2/Y BUFX2_99/A NAND3X1_7/B DFFSR_92/S NAND3X1
XFILL_20_DFFPOSX1_44 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_19_DFFSR_159 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_33_DFFSR_263 OR2X2_1/gnd DFFSR_51/S FILL
XNOR2X1_41 NOR2X1_41/A NOR2X1_41/B DFFSR_1/gnd NOR2X1_41/Y DFFSR_81/S NOR2X1
XFILL_4_NAND3X1_3 BUFX2_99/A DFFSR_92/S FILL
XFILL_23_DFFSR_266 INVX1_67/gnd DFFSR_201/S FILL
XFILL_4_NAND3X1_247 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_4_NOR2X1_38 INVX1_3/gnd DFFSR_79/S FILL
XFILL_13_DFFSR_269 INVX1_67/gnd DFFSR_201/S FILL
XFILL_12_CLKBUF1_11 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_7_OAI21X1_103 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_7_DFFSR_58 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_35_DFFSR_11 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_13_DFFSR_91 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_24_DFFSR_51 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_11_CLKBUF1_14 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_5_DFFSR_156 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_10_CLKBUF1_17 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_46_DFFSR_187 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_5_NAND3X1_181 INVX1_39/gnd DFFSR_54/S FILL
XFILL_9_DFFSR_263 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_36_DFFSR_190 INVX1_39/gnd DFFSR_34/S FILL
XFILL_26_DFFSR_193 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_9_CLKBUF1_20 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_7_DFFSR_5 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_16_DFFSR_196 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_8_CLKBUF1_23 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_6_NAND3X1_115 BUFX2_79/A DFFSR_7/S FILL
XFILL_7_CLKBUF1_26 INVX1_1/gnd DFFSR_53/S FILL
XFILL_10_DFFPOSX1_19 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_32_DFFSR_58 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_4_INVX1_52 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_21_DFFSR_98 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_43_DFFSR_18 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_6_CLKBUF1_29 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_1_NOR2X1_75 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_49_DFFSR_114 NOR3X1_6/gnd DFFSR_91/S FILL
XNAND3X1_151 AOI21X1_14/A AOI21X1_12/C AOI21X1_14/B DFFSR_1/gnd NAND3X1_152/B DFFSR_81/S
+ NAND3X1
XFILL_5_CLKBUF1_32 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_39_DFFSR_117 BUFX2_77/gnd DFFSR_98/S FILL
XCLKBUF1_29 BUFX2_6/Y XOR2X1_4/gnd CLKBUF1_29/Y DFFSR_91/S CLKBUF1
XFILL_4_CLKBUF1_35 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_2_DFFSR_193 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_3_BUFX2_43 AND2X2_38/B DFFSR_23/S FILL
XFILL_5_OR2X2_5 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_29_DFFSR_120 INVX1_3/gnd DFFSR_23/S FILL
XFILL_43_DFFSR_224 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_3_CLKBUF1_38 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_8_AND2X2_34 AND2X2_38/B DFFSR_59/S FILL
XFILL_19_DFFSR_123 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_33_DFFSR_227 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_2_CLKBUF1_41 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_31_DFFSR_9 BUFX2_79/A DFFSR_6/S FILL
XFILL_23_DFFSR_230 INVX1_67/gnd DFFSR_201/S FILL
XFILL_4_NAND3X1_211 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_1_CLKBUF1_44 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_1_INVX1_99 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_40_DFFSR_65 BUFX2_79/A DFFSR_7/S FILL
XFILL_13_DFFSR_233 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_0_DFFPOSX1_30 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_0_CLKBUF1_47 BUFX2_98/A DFFSR_32/S FILL
XFILL_16_2 INVX1_39/gnd DFFSR_34/S FILL
XFILL_7_DFFSR_22 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_24_DFFSR_15 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_13_DFFSR_55 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_5_DFFSR_120 INVX1_3/gnd DFFSR_23/S FILL
XFILL_0_BUFX2_90 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_46_DFFSR_151 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_5_NAND3X1_145 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_9_DFFSR_227 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_31_2_0 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_36_DFFSR_154 BUFX2_99/A DFFSR_7/S FILL
XFILL_50_DFFSR_258 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_6_NOR2X1_3 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_26_DFFSR_157 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_40_DFFSR_261 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_2_INVX1_204 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_48_DFFSR_72 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_29_4_1 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_16_DFFSR_160 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_30_DFFSR_264 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_1_NAND3X1_4 BUFX2_79/A DFFSR_7/S FILL
XFILL_20_DFFSR_267 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_32_DFFSR_22 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_4_DFFSR_69 BUFX2_98/A DFFSR_32/S FILL
XFILL_21_DFFSR_62 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_27_6_2 INVX1_3/gnd DFFSR_79/S FILL
XFILL_19_DFFPOSX1_38 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_1_NOR2X1_39 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_10_DFFSR_270 INVX1_39/gnd DFFSR_54/S FILL
XNAND3X1_115 BUFX2_96/A AND2X2_16/Y BUFX2_33/Y BUFX2_79/A AND2X2_25/A DFFSR_7/S NAND3X1
XFILL_9_5_1 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_3_NAND3X1_241 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_2_DFFSR_157 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_43_DFFSR_188 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_6_DFFSR_264 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_33_DFFSR_191 INVX1_67/gnd DFFSR_175/S FILL
XFILL_4_NAND3X1_175 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_23_DFFSR_194 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_40_DFFSR_29 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_1_INVX1_63 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_29_DFFSR_69 BUFX2_98/A DFFSR_32/S FILL
XFILL_13_DFFSR_197 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_0_CLKBUF1_11 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_9_DFFPOSX1_49 BUFX2_99/A DFFSR_92/S FILL
XFILL_13_DFFSR_19 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_0_BUFX2_54 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_5_NAND3X1_109 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_46_DFFSR_115 INVX1_1/gnd DFFSR_97/S FILL
XFILL_9_DFFSR_191 INVX1_67/gnd DFFSR_175/S FILL
XFILL_36_DFFSR_118 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_50_DFFSR_222 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_18_DFFSR_3 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_26_DFFSR_121 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_40_DFFSR_225 INVX1_67/gnd DFFSR_175/S FILL
XFILL_48_DFFSR_36 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_37_DFFSR_76 BUFX2_79/A DFFSR_7/S FILL
XFILL_2_INVX1_168 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_5_AND2X2_35 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_16_DFFSR_124 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_30_DFFSR_228 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_37_1_2 BUFX2_99/A DFFSR_7/S FILL
XFILL_6_AOI21X1_3 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_20_DFFSR_231 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_4_DFFSR_33 BUFX2_98/A DFFSR_32/S FILL
XFILL_21_DFFSR_26 BUFX2_79/A DFFSR_6/S FILL
XFILL_10_DFFSR_66 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_2_BUFX2_4 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_10_DFFSR_234 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_3_NAND3X1_205 INVX1_1/gnd DFFSR_53/S FILL
XFILL_2_DFFSR_121 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_43_DFFSR_152 INVX1_1/gnd DFFSR_53/S FILL
XFILL_45_DFFSR_83 INVX1_3/gnd DFFSR_79/S FILL
XFILL_6_DFFSR_228 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_33_DFFSR_155 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_47_DFFSR_259 BUFX2_79/A DFFSR_6/S FILL
XFILL_23_DFFSR_158 INVX1_3/gnd DFFSR_23/S FILL
XFILL_4_NAND3X1_139 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_37_DFFSR_262 BUFX2_98/A DFFSR_32/S FILL
XFILL_1_INVX1_27 BUFX2_99/A DFFSR_7/S FILL
XFILL_1_DFFSR_80 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_29_DFFSR_33 BUFX2_98/A DFFSR_32/S FILL
XFILL_18_DFFSR_73 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_8_NAND3X1_2 BUFX2_99/A DFFSR_7/S FILL
XFILL_13_DFFSR_161 INVX1_67/gnd DFFSR_175/S FILL
XFILL_27_DFFSR_265 INVX1_67/gnd DFFSR_175/S FILL
XFILL_9_DFFPOSX1_13 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_23_DFFPOSX1_2 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_6_NAND2X1_175 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_17_DFFSR_268 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_22_DFFPOSX1_5 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_0_BUFX2_18 BUFX2_98/A DFFSR_32/S FILL
XFILL_21_DFFPOSX1_8 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_9_DFFSR_155 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_18_DFFPOSX1_32 INVX1_67/gnd DFFSR_201/S FILL
XFILL_50_DFFSR_186 BUFX2_99/A DFFSR_92/S FILL
XFILL_40_DFFSR_189 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_37_DFFSR_40 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_9_DFFSR_87 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_2_INVX1_132 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_26_DFFSR_80 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_2_NAND3X1_235 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_3_DFFSR_265 INVX1_67/gnd DFFSR_175/S FILL
XFILL_30_DFFSR_192 INVX1_1/gnd DFFSR_97/S FILL
XFILL_20_DFFSR_195 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_10_DFFSR_30 BUFX2_98/A DFFSR_32/S FILL
XFILL_10_DFFSR_198 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_5_NOR2X1_74 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_3_NAND3X1_169 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_18_NOR3X1_4 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_8_DFFPOSX1_43 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_43_DFFSR_116 INVX1_3/gnd DFFSR_23/S FILL
XFILL_34_DFFSR_87 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_45_DFFSR_47 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_6_DFFSR_192 INVX1_1/gnd DFFSR_97/S FILL
XFILL_33_DFFSR_119 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_47_DFFSR_223 INVX1_39/gnd DFFSR_34/S FILL
XFILL_23_DFFSR_122 BUFX2_79/A DFFSR_7/S FILL
XFILL_4_NAND3X1_103 AND2X2_38/B DFFSR_23/S FILL
XFILL_37_DFFSR_226 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_1_DFFSR_44 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_18_DFFSR_37 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_2_AND2X2_36 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_5_BUFX2_72 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_13_DFFSR_125 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_27_DFFSR_229 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_3_AOI21X1_4 BUFX2_98/A DFFSR_32/S FILL
XFILL_6_NAND2X1_139 INVX1_1/gnd DFFSR_97/S FILL
XFILL_17_DFFSR_232 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_6_DFFSR_2 BUFX2_79/A DFFSR_7/S FILL
XFILL_11_XOR2X1_7 BUFX2_98/A DFFSR_6/S FILL
XFILL_9_DFFSR_119 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_42_DFFSR_94 BUFX2_77/gnd DFFSR_98/S FILL
XNAND2X1_175 AOI21X1_66/Y AOI21X1_68/A XOR2X1_4/gnd AOI21X1_67/A DFFSR_91/S NAND2X1
XFILL_50_DFFSR_150 AND2X2_38/B DFFSR_23/S FILL
XFILL_8_AOI21X1_67 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_40_DFFSR_153 INVX1_67/gnd DFFSR_201/S FILL
XFILL_3_AND2X2_3 INVX1_1/gnd DFFSR_53/S FILL
XFILL_26_DFFSR_44 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_7_AOI21X1_70 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_9_DFFSR_51 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_15_DFFSR_84 BUFX2_99/A DFFSR_7/S FILL
XFILL_2_NAND3X1_199 INVX1_1/gnd DFFSR_97/S FILL
XFILL_3_DFFSR_229 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_30_DFFSR_156 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_44_DFFSR_260 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_4_OR2X2_2 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_20_DFFSR_159 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_34_DFFSR_263 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_5_NAND3X1_3 BUFX2_99/A DFFSR_92/S FILL
XFILL_10_DFFSR_162 BUFX2_99/A DFFSR_92/S FILL
XFILL_24_DFFSR_266 INVX1_67/gnd DFFSR_201/S FILL
XFILL_30_DFFSR_6 BUFX2_79/A DFFSR_6/S FILL
XFILL_5_NOR2X1_38 INVX1_3/gnd DFFSR_79/S FILL
XFILL_3_NAND3X1_133 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_14_DFFSR_269 INVX1_67/gnd DFFSR_201/S FILL
XFILL_38_2_0 BUFX2_79/A DFFSR_7/S FILL
XFILL_5_NAND2X1_169 INVX1_1/gnd DFFSR_53/S FILL
XFILL_6_DFFSR_98 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_23_DFFSR_91 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_34_DFFSR_51 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_45_DFFSR_11 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_6_DFFSR_156 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_36_4_1 BUFX2_99/A DFFSR_92/S FILL
XFILL_47_DFFSR_187 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_11_DFFPOSX1_2 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_37_DFFSR_190 INVX1_39/gnd DFFSR_34/S FILL
XBUFX2_76 BUFX2_76/A OR2X2_2/gnd dout[5] DFFSR_216/S BUFX2
XFILL_0_DFFSR_266 INVX1_67/gnd DFFSR_201/S FILL
XFILL_5_BUFX2_36 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_10_DFFPOSX1_5 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_34_6_2 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_17_DFFPOSX1_26 AND2X2_38/B DFFSR_23/S FILL
XFILL_27_DFFSR_193 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_6_NAND2X1_103 AND2X2_38/B DFFSR_23/S FILL
XFILL_17_DFFSR_196 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_1_NAND3X1_229 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_9_DFFPOSX1_8 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_42_DFFSR_58 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_3_INVX1_92 AND2X2_38/B DFFSR_23/S FILL
XFILL_31_DFFSR_98 BUFX2_77/gnd DFFSR_98/S FILL
XNAND2X1_139 DFFSR_91/S DFFSR_272/Q INVX1_1/gnd NAND2X1_139/Y DFFSR_97/S NAND2X1
XFILL_2_NOR2X1_75 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_50_DFFSR_114 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_8_AOI21X1_31 INVX1_39/gnd DFFSR_34/S FILL
XFILL_27_DFFPOSX1_15 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_40_DFFSR_117 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_9_DFFSR_15 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_7_AOI21X1_34 INVX1_39/gnd DFFSR_34/S FILL
XFILL_15_DFFSR_48 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_2_NAND3X1_163 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_3_DFFSR_193 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_2_BUFX2_83 BUFX2_79/A DFFSR_7/S FILL
XFILL_30_DFFSR_120 INVX1_3/gnd DFFSR_23/S FILL
XFILL_6_AOI21X1_37 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_44_DFFSR_224 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_9_AND2X2_34 AND2X2_38/B DFFSR_59/S FILL
XFILL_7_DFFPOSX1_37 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_20_DFFSR_123 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_34_DFFSR_227 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_5_AOI21X1_40 INVX1_39/gnd DFFSR_54/S FILL
XAOI21X1_37 AOI21X1_37/A AOI21X1_37/B XOR2X1_6/Y OR2X2_3/gnd OAI21X1_80/B DFFSR_4/S
+ AOI21X1
XFILL_10_DFFSR_126 BUFX2_99/A DFFSR_7/S FILL
XFILL_4_AOI21X1_43 INVX1_3/gnd DFFSR_79/S FILL
XFILL_24_DFFSR_230 INVX1_67/gnd DFFSR_201/S FILL
XFILL_0_AOI21X1_5 INVX1_3/gnd DFFSR_23/S FILL
XFILL_50_DFFSR_65 BUFX2_79/A DFFSR_7/S FILL
XFILL_3_AOI21X1_46 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_14_DFFSR_233 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_2_AOI21X1_49 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_5_NAND2X1_133 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_34_DFFSR_15 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_23_DFFSR_55 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_12_DFFSR_95 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_6_DFFSR_62 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_1_AOI21X1_52 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_6_DFFSR_120 INVX1_3/gnd DFFSR_23/S FILL
XFILL_47_DFFSR_151 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_0_AOI21X1_55 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_44_1_2 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_37_DFFSR_154 BUFX2_99/A DFFSR_7/S FILL
XFILL_51_DFFSR_258 DFFSR_5/gnd DFFSR_5/S FILL
XBUFX2_40 rst INVX1_1/gnd BUFX2_40/Y DFFSR_97/S BUFX2
XFILL_0_DFFSR_230 INVX1_67/gnd DFFSR_201/S FILL
XFILL_27_DFFSR_157 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_3_OAI21X1_115 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_41_DFFSR_261 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_26_DFFPOSX1_45 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_3_INVX1_204 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_17_DFFSR_160 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_8_OAI21X1_79 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_31_DFFSR_264 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_1_NAND3X1_193 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_2_NAND3X1_4 BUFX2_79/A DFFSR_7/S FILL
XFILL_7_OAI21X1_82 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_21_DFFSR_267 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_42_DFFSR_22 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_3_INVX1_56 BUFX2_98/A DFFSR_6/S FILL
XFILL_31_DFFSR_62 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_2_NOR2X1_39 OR2X2_6/gnd DFFSR_92/S FILL
XNAND2X1_103 OAI21X1_69/Y NAND3X1_214/B AND2X2_38/B INVX1_179/A DFFSR_23/S NAND2X1
XFILL_11_DFFSR_270 INVX1_39/gnd DFFSR_54/S FILL
XFILL_6_OAI21X1_85 INVX1_39/gnd DFFSR_54/S FILL
XFILL_5_OAI21X1_88 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_12_0_0 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_1_BUFX2_1 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_15_DFFSR_12 DFFSR_8/gnd DFFSR_8/S FILL
XOAI21X1_85 DFFSR_54/S INVX1_181/Y OAI21X1_85/C INVX1_39/gnd DFFSR_257/D DFFSR_54/S
+ OAI21X1
XFILL_2_NAND3X1_127 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_3_DFFSR_157 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_4_OAI21X1_91 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_2_BUFX2_47 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_44_DFFSR_188 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_3_OAI21X1_94 INVX1_67/gnd DFFSR_175/S FILL
XFILL_10_2_1 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_7_DFFSR_264 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_4_NAND2X1_163 INVX1_67/gnd DFFSR_201/S FILL
XFILL_34_DFFSR_191 INVX1_67/gnd DFFSR_175/S FILL
XFILL_2_OAI21X1_97 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_24_DFFSR_194 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_50_DFFSR_29 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_39_DFFSR_69 BUFX2_98/A DFFSR_32/S FILL
XFILL_3_AOI21X1_10 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_14_DFFSR_197 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_3_3 INVX1_67/gnd DFFSR_201/S FILL
XFILL_2_AOI21X1_13 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_16_DFFPOSX1_20 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_23_DFFSR_19 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_6_DFFSR_26 BUFX2_79/A DFFSR_6/S FILL
XFILL_12_DFFSR_59 AND2X2_38/B DFFSR_59/S FILL
XFILL_1_AOI21X1_16 INVX1_67/gnd DFFSR_175/S FILL
XFILL_47_DFFSR_115 INVX1_1/gnd DFFSR_97/S FILL
XFILL_0_NAND3X1_223 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_0_AOI21X1_19 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_37_DFFSR_118 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_5_NOR2X1_7 BUFX2_98/A DFFSR_32/S FILL
XFILL_0_DFFSR_194 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_27_DFFSR_121 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_42_DFFSR_9 BUFX2_79/A DFFSR_6/S FILL
XFILL_41_DFFSR_225 INVX1_67/gnd DFFSR_175/S FILL
XFILL_47_DFFSR_76 BUFX2_79/A DFFSR_7/S FILL
XFILL_3_INVX1_168 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_6_AND2X2_35 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_17_DFFSR_124 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_8_OAI21X1_43 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_1_NAND3X1_157 INVX1_3/gnd DFFSR_23/S FILL
XFILL_31_DFFSR_228 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_7_AOI21X1_3 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_7_OAI21X1_46 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_6_NAND2X1_64 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_21_DFFSR_231 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_3_INVX1_20 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_3_DFFSR_73 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_20_DFFSR_66 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_31_DFFSR_26 BUFX2_79/A DFFSR_6/S FILL
XFILL_6_DFFPOSX1_31 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_11_DFFSR_234 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_5_NAND2X1_67 AND2X2_38/B DFFSR_59/S FILL
XFILL_6_OAI21X1_49 DFFSR_34/gnd DFFSR_1/S FILL
XNAND2X1_64 NAND2X1_64/A NAND2X1_64/B DFFSR_46/gnd OAI21X1_25/C DFFSR_62/S NAND2X1
XFILL_4_NAND2X1_70 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_5_OAI21X1_52 XOR2X1_1/gnd DFFSR_208/S FILL
XOAI21X1_49 INVX1_145/Y INVX1_159/Y AND2X2_35/Y DFFSR_34/gnd OAI21X1_49/Y DFFSR_1/S
+ OAI21X1
XFILL_3_DFFSR_121 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_3_NAND2X1_73 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_4_OAI21X1_55 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_2_BUFX2_11 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_7_XOR2X1_3 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_44_DFFSR_152 INVX1_1/gnd DFFSR_53/S FILL
XFILL_15_DFFPOSX1_50 INVX1_1/gnd DFFSR_53/S FILL
XFILL_2_NAND2X1_76 INVX1_3/gnd DFFSR_23/S FILL
XFILL_3_OAI21X1_58 INVX1_39/gnd DFFSR_54/S FILL
XFILL_7_DFFSR_228 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_34_DFFSR_155 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_4_NAND2X1_127 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_48_DFFSR_259 BUFX2_79/A DFFSR_6/S FILL
XFILL_2_OAI21X1_61 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_1_NAND2X1_79 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_11_AOI22X1_27 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_24_DFFSR_158 INVX1_3/gnd DFFSR_23/S FILL
XFILL_1_OAI21X1_64 INVX1_1/gnd DFFSR_53/S FILL
XFILL_0_NAND2X1_82 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_0_INVX1_67 INVX1_67/gnd DFFSR_201/S FILL
XFILL_38_DFFSR_262 BUFX2_98/A DFFSR_32/S FILL
XFILL_39_DFFSR_33 BUFX2_98/A DFFSR_32/S FILL
XFILL_0_INVX1_205 BUFX2_99/A DFFSR_92/S FILL
XFILL_28_DFFSR_73 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_14_DFFSR_161 INVX1_67/gnd DFFSR_175/S FILL
XFILL_0_OAI21X1_67 INVX1_1/gnd DFFSR_97/S FILL
XFILL_28_DFFSR_265 INVX1_67/gnd DFFSR_175/S FILL
XFILL_2_OAI21X1_109 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_25_DFFPOSX1_39 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_18_DFFSR_268 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_12_DFFSR_23 AND2X2_38/B DFFSR_23/S FILL
XFILL_0_NAND3X1_187 BUFX2_7/gnd DFFSR_216/S FILL
XDFFSR_3 DFFSR_3/Q DFFSR_3/CLK DFFSR_3/R DFFSR_3/S DFFSR_3/D OR2X2_4/gnd DFFSR_3/S
+ DFFSR
XFILL_3_NOR3X1_4 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_0_DFFSR_158 INVX1_3/gnd DFFSR_23/S FILL
XDFFSR_268 INVX1_193/A CLKBUF1_48/Y DFFSR_266/R DFFSR_51/S DFFSR_268/D OR2X2_1/gnd
+ DFFSR_51/S DFFSR
XFILL_41_DFFSR_189 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_47_DFFSR_40 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_3_INVX1_132 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_36_DFFSR_80 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_4_DFFSR_265 INVX1_67/gnd DFFSR_175/S FILL
XFILL_1_NAND3X1_121 INVX1_1/gnd DFFSR_97/S FILL
XFILL_31_DFFSR_192 INVX1_1/gnd DFFSR_97/S FILL
XFILL_45_2_0 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_7_OAI21X1_10 BUFX2_79/A DFFSR_7/S FILL
XFILL_6_NAND2X1_28 AND2X2_38/B DFFSR_59/S FILL
XFILL_21_DFFSR_195 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_3_DFFSR_37 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_20_DFFSR_30 BUFX2_98/A DFFSR_32/S FILL
XFILL_5_NAND2X1_31 INVX1_3/gnd DFFSR_23/S FILL
XFILL_11_DFFSR_198 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_3_NAND2X1_157 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_6_OAI21X1_13 INVX1_39/gnd DFFSR_54/S FILL
XNAND2X1_28 NOR2X1_30/Y BUFX2_25/Y AND2X2_38/B OAI22X1_43/B DFFSR_59/S NAND2X1
XFILL_43_4_1 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_5_OAI21X1_16 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_4_NAND2X1_34 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_6_NOR2X1_74 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_8_8 BUFX2_7/gnd DFFSR_151/S FILL
XOAI21X1_13 INVX1_96/Y OAI21X1_9/B OAI21X1_13/C INVX1_39/gnd NOR2X1_48/B DFFSR_54/S
+ OAI21X1
XFILL_3_NAND2X1_37 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_4_OAI21X1_19 BUFX2_98/A DFFSR_32/S FILL
XDFFPOSX1_31 NAND2X1_151/B CLKBUF1_45/Y AOI21X1_52/Y XOR2X1_4/gnd DFFSR_97/S DFFPOSX1
XFILL_44_DFFSR_116 INVX1_3/gnd DFFSR_23/S FILL
XFILL_29_DFFSR_3 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_41_6_2 BUFX2_98/A DFFSR_32/S FILL
XFILL_2_NAND2X1_40 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_3_OAI21X1_22 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_15_DFFPOSX1_14 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_44_DFFSR_87 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_7_DFFSR_192 INVX1_1/gnd DFFSR_97/S FILL
XFILL_34_DFFSR_119 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_1_NAND2X1_43 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_48_DFFSR_223 INVX1_39/gnd DFFSR_34/S FILL
XFILL_2_OAI21X1_25 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_24_DFFSR_122 BUFX2_79/A DFFSR_7/S FILL
XFILL_8_NAND3X1_99 OR2X2_1/gnd DFFSR_51/S FILL
XAOI21X1_7 AOI21X1_7/A AOI21X1_7/B AOI21X1_7/C OR2X2_2/gnd INVX1_153/A DFFSR_175/S
+ AOI21X1
XFILL_1_OAI21X1_28 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_0_NAND2X1_46 INVX1_39/gnd DFFSR_34/S FILL
XFILL_28_DFFSR_37 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_38_DFFSR_226 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_0_DFFSR_84 BUFX2_99/A DFFSR_7/S FILL
XFILL_0_INVX1_31 INVX1_1/gnd DFFSR_53/S FILL
XFILL_0_INVX1_169 INVX1_39/gnd DFFSR_34/S FILL
XFILL_17_DFFSR_77 BUFX2_98/A DFFSR_32/S FILL
XFILL_3_AND2X2_36 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_14_DFFSR_125 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_0_OAI21X1_31 AND2X2_38/B DFFSR_23/S FILL
XFILL_28_DFFSR_229 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_4_AOI21X1_4 BUFX2_98/A DFFSR_32/S FILL
XFILL_18_DFFSR_232 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_0_NAND3X1_151 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_5_DFFPOSX1_25 BUFX2_79/A DFFSR_6/S FILL
XFILL_0_DFFSR_122 BUFX2_79/A DFFSR_7/S FILL
XDFFSR_232 DFFSR_232/Q CLKBUF1_14/Y BUFX2_64/Y DFFSR_54/S DFFSR_224/Q DFFSR_46/gnd
+ DFFSR_54/S DFFSR
XFILL_41_DFFSR_153 INVX1_67/gnd DFFSR_201/S FILL
XFILL_8_DFFSR_91 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_36_DFFSR_44 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_25_DFFSR_84 BUFX2_99/A DFFSR_7/S FILL
XFILL_4_DFFSR_229 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_31_DFFSR_156 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_45_DFFSR_260 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_4_AOI22X1_12 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_21_DFFSR_159 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_14_DFFPOSX1_44 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_35_DFFSR_263 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_3_AOI22X1_15 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_6_NAND3X1_3 BUFX2_99/A DFFSR_92/S FILL
XFILL_3_NAND2X1_121 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_11_DFFSR_162 BUFX2_99/A DFFSR_92/S FILL
XFILL_25_DFFSR_266 INVX1_67/gnd DFFSR_201/S FILL
XFILL_2_AOI22X1_18 OR2X2_1/gnd DFFSR_59/S FILL
XINVX1_5 INVX1_5/A BUFX2_8/gnd INVX1_5/Y DFFSR_81/S INVX1
XFILL_6_NOR2X1_38 INVX1_3/gnd DFFSR_79/S FILL
XFILL_15_DFFSR_269 INVX1_67/gnd DFFSR_201/S FILL
XFILL_51_1_2 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_1_AOI22X1_21 AND2X2_38/B DFFSR_59/S FILL
XFILL_10_OAI22X1_42 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_0_AOI22X1_24 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_1_OAI21X1_103 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_33_DFFSR_91 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_44_DFFSR_51 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_7_DFFSR_156 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_24_DFFPOSX1_33 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_48_DFFSR_187 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_9_OAI22X1_45 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_8_NAND3X1_63 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_0_NAND2X1_10 BUFX2_79/A DFFSR_7/S FILL
XFILL_38_DFFSR_190 INVX1_39/gnd DFFSR_34/S FILL
XFILL_0_DFFSR_48 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_8_NAND3X1_236 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_17_DFFSR_41 BUFX2_98/A DFFSR_6/S FILL
XFILL_0_INVX1_133 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_1_DFFSR_266 INVX1_67/gnd DFFSR_201/S FILL
XFILL_7_NAND3X1_66 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_8_OAI22X1_48 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_4_BUFX2_76 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_28_DFFSR_193 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_6_NAND3X1_69 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_7_OAI22X1_51 INVX1_39/gnd DFFSR_54/S FILL
XFILL_18_DFFSR_196 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_19_0_0 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_5_NAND3X1_72 INVX1_39/gnd DFFSR_34/S FILL
XNAND3X1_69 DFFSR_193/D BUFX2_31/Y BUFX2_24/Y BUFX2_7/gnd NAND3X1_71/A DFFSR_216/S
+ NAND3X1
XFILL_0_NAND3X1_115 BUFX2_79/A DFFSR_7/S FILL
XFILL_4_NAND3X1_75 BUFX2_79/A DFFSR_7/S FILL
XFILL_41_DFFSR_98 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_3_NOR2X1_75 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_17_2_1 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_51_DFFSR_114 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_3_NAND3X1_78 NOR3X1_6/gnd DFFSR_79/S FILL
XDFFSR_196 DFFSR_204/D CLKBUF1_21/Y BUFX2_68/Y DFFSR_151/S DFFSR_196/D XOR2X1_1/gnd
+ DFFSR_151/S DFFSR
XFILL_2_NAND2X1_151 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_41_DFFSR_117 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_2_AND2X2_7 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_8_DFFSR_55 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_2_NAND3X1_81 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_25_DFFSR_48 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_14_DFFSR_88 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_4_DFFSR_193 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_31_DFFSR_120 INVX1_3/gnd DFFSR_23/S FILL
XFILL_15_4_2 INVX1_39/gnd DFFSR_34/S FILL
XFILL_1_NAND3X1_84 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_45_DFFSR_224 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_21_DFFSR_123 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_0_NAND3X1_87 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_35_DFFSR_227 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_0_AND2X2_37 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_11_DFFSR_126 BUFX2_99/A DFFSR_7/S FILL
XFILL_25_DFFSR_230 INVX1_67/gnd DFFSR_201/S FILL
XFILL_1_AOI21X1_5 INVX1_3/gnd DFFSR_23/S FILL
XFILL_15_DFFSR_233 OR2X2_2/gnd DFFSR_175/S FILL
XINVX1_89 INVX1_89/A OR2X2_1/gnd INVX1_89/Y DFFSR_51/S INVX1
XFILL_44_DFFSR_15 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_33_DFFSR_55 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_22_DFFSR_95 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_7_DFFSR_120 INVX1_3/gnd DFFSR_23/S FILL
XFILL_9_NAND3X1_24 INVX1_1/gnd DFFSR_97/S FILL
XFILL_48_DFFSR_151 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_8_NAND3X1_27 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_38_DFFSR_154 BUFX2_99/A DFFSR_7/S FILL
XFILL_0_DFFSR_12 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_8_NAND3X1_200 OR2X2_6/gnd DFFSR_53/S FILL
XINVX1_207 BUFX2_35/Y DFFSR_1/gnd DFFSR_274/R DFFSR_1/S INVX1
XFILL_1_DFFSR_230 INVX1_67/gnd DFFSR_201/S FILL
XFILL_8_OAI22X1_12 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_7_NAND3X1_30 BUFX2_79/A DFFSR_6/S FILL
XFILL_4_BUFX2_40 INVX1_1/gnd DFFSR_97/S FILL
XFILL_28_DFFSR_157 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_4_DFFPOSX1_19 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_1_NAND2X1_181 BUFX2_99/A DFFSR_92/S FILL
XFILL_4_INVX1_204 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_6_NAND3X1_33 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_42_DFFSR_261 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_7_OAI22X1_15 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_18_DFFSR_160 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_32_DFFSR_264 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_6_OAI22X1_18 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_5_NAND3X1_36 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_41_DFFSR_6 BUFX2_79/A DFFSR_6/S FILL
XFILL_3_NAND3X1_4 BUFX2_79/A DFFSR_7/S FILL
XNAND3X1_33 DFFSR_61/D BUFX2_15/Y BUFX2_14/Y DFFSR_8/gnd NAND3X1_33/Y DFFSR_8/S NAND3X1
XFILL_22_DFFSR_267 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_4_NAND3X1_39 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_5_OAI22X1_21 BUFX2_98/A DFFSR_32/S FILL
XFILL_2_INVX1_96 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_41_DFFSR_62 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_3_NOR2X1_39 OR2X2_6/gnd DFFSR_92/S FILL
XOAI22X1_18 INVX1_42/Y OAI22X1_6/B INVX1_43/Y OAI22X1_6/D OR2X2_4/gnd NOR2X1_22/A
+ DFFSR_3/S OAI22X1
XFILL_13_DFFPOSX1_38 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_12_DFFSR_270 INVX1_39/gnd DFFSR_54/S FILL
XFILL_4_OAI22X1_24 BUFX2_98/A DFFSR_32/S FILL
XFILL_3_NAND3X1_42 BUFX2_79/A DFFSR_6/S FILL
XFILL_2_NAND2X1_115 DFFSR_28/gnd DFFSR_3/S FILL
XDFFSR_160 DFFSR_160/Q CLKBUF1_39/Y BUFX2_63/Y DFFSR_97/S DFFSR_136/Q XOR2X1_4/gnd
+ DFFSR_97/S DFFSR
XFILL_3_OAI22X1_27 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_8_DFFSR_19 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_2_NAND3X1_45 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_25_DFFSR_12 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_14_DFFSR_52 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_4_DFFSR_157 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_1_BUFX2_87 INVX1_1/gnd DFFSR_53/S FILL
XFILL_1_NAND3X1_48 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_2_OAI22X1_30 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_45_DFFSR_188 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_8_DFFSR_264 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_0_NAND3X1_51 BUFX2_99/A DFFSR_7/S FILL
XFILL_1_OAI22X1_33 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_35_DFFSR_191 INVX1_67/gnd DFFSR_175/S FILL
XFILL_5_0_2 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_23_DFFPOSX1_27 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_0_OAI22X1_36 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_25_DFFSR_194 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_49_DFFSR_69 BUFX2_98/A DFFSR_32/S FILL
XFILL_7_NAND3X1_230 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_15_DFFSR_197 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_3_DFFPOSX1_49 BUFX2_99/A DFFSR_92/S FILL
XINVX1_53 DFFSR_56/D DFFSR_8/gnd INVX1_53/Y DFFSR_60/S INVX1
XFILL_33_DFFSR_19 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_5_DFFSR_66 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_11_DFFSR_99 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_22_DFFSR_59 AND2X2_38/B DFFSR_59/S FILL
XFILL_0_NOR2X1_76 INVX1_3/gnd DFFSR_79/S FILL
XFILL_48_DFFSR_115 INVX1_1/gnd DFFSR_97/S FILL
XFILL_38_DFFSR_118 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_52_2_0 BUFX2_77/gnd DFFSR_98/S FILL
XINVX1_171 XOR2X1_8/A BUFX2_98/A INVX1_171/Y DFFSR_6/S INVX1
XFILL_8_NAND3X1_164 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_1_DFFSR_194 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_28_DFFSR_121 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_1_NAND2X1_145 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_42_DFFSR_225 INVX1_67/gnd DFFSR_175/S FILL
XFILL_4_INVX1_168 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_7_AND2X2_35 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_50_4_1 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_18_DFFSR_124 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_32_DFFSR_228 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_8_AOI21X1_3 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_22_DFFSR_231 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_30_DFFSR_66 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_41_DFFSR_26 BUFX2_79/A DFFSR_6/S FILL
XFILL_2_INVX1_60 INVX1_39/gnd DFFSR_34/S FILL
XFILL_48_6_2 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_12_DFFSR_234 OR2X2_3/gnd DFFSR_4/S FILL
XDFFSR_124 BUFX2_85/A CLKBUF1_8/Y DFFSR_1/R DFFSR_59/S INVX1_30/A OR2X2_1/gnd DFFSR_59/S
+ DFFSR
XFILL_14_DFFSR_16 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_4_DFFSR_121 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_1_BUFX2_51 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_1_NAND3X1_12 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_45_DFFSR_152 INVX1_1/gnd DFFSR_53/S FILL
XFILL_0_NAND3X1_15 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_8_DFFSR_228 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_8_DFFSR_9 BUFX2_79/A DFFSR_6/S FILL
XFILL_35_DFFSR_155 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_49_DFFSR_259 BUFX2_79/A DFFSR_6/S FILL
XFILL_9_OAI21X1_116 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_25_DFFSR_158 INVX1_3/gnd DFFSR_23/S FILL
XFILL_39_DFFSR_262 BUFX2_98/A DFFSR_32/S FILL
XFILL_49_DFFSR_33 BUFX2_98/A DFFSR_32/S FILL
XFILL_1_INVX1_205 BUFX2_99/A DFFSR_92/S FILL
XFILL_38_DFFSR_73 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_15_DFFSR_161 INVX1_67/gnd DFFSR_175/S FILL
XFILL_16_5_0 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_7_NAND3X1_194 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_29_DFFSR_265 INVX1_67/gnd DFFSR_175/S FILL
XFILL_0_NAND3X1_5 BUFX2_99/A DFFSR_7/S FILL
XFILL_3_DFFPOSX1_13 BUFX2_8/gnd DFFSR_81/S FILL
XDFFSR_70 DFFSR_70/Q CLKBUF1_5/Y DFFSR_9/R DFFSR_8/S DFFSR_14/Q DFFSR_28/gnd DFFSR_8/S
+ DFFSR
XFILL_0_NAND2X1_175 XOR2X1_4/gnd DFFSR_91/S FILL
XINVX1_17 DFFSR_11/D AND2X2_38/B INVX1_17/Y DFFSR_59/S INVX1
XFILL_19_DFFSR_268 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_5_DFFSR_30 BUFX2_98/A DFFSR_32/S FILL
XFILL_11_DFFSR_63 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_22_DFFSR_23 AND2X2_38/B DFFSR_23/S FILL
XFILL_0_NOR2X1_40 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_8_NAND3X1_128 NOR3X1_6/gnd DFFSR_79/S FILL
XINVX1_135 INVX1_135/A BUFX2_8/gnd INVX1_135/Y DFFSR_51/S INVX1
XFILL_1_DFFSR_158 INVX1_3/gnd DFFSR_23/S FILL
XFILL_12_DFFPOSX1_32 INVX1_67/gnd DFFSR_201/S FILL
XFILL_1_NAND2X1_109 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_42_DFFSR_189 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_46_DFFSR_80 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_5_DFFSR_265 INVX1_67/gnd DFFSR_175/S FILL
XFILL_32_DFFSR_192 INVX1_1/gnd DFFSR_97/S FILL
XFILL_22_DFFSR_195 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_19_DFFSR_70 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_2_INVX1_24 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_30_DFFSR_30 BUFX2_98/A DFFSR_32/S FILL
XFILL_2_DFFSR_77 BUFX2_98/A DFFSR_32/S FILL
XFILL_12_DFFSR_198 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_22_DFFPOSX1_21 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_1_BUFX2_15 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_6_NAND3X1_224 INVX1_39/gnd DFFSR_54/S FILL
XFILL_6_XOR2X1_7 BUFX2_98/A DFFSR_6/S FILL
XFILL_45_DFFSR_116 INVX1_3/gnd DFFSR_23/S FILL
XFILL_2_DFFPOSX1_43 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_8_DFFSR_192 INVX1_1/gnd DFFSR_97/S FILL
XFILL_35_DFFSR_119 OR2X2_4/gnd DFFSR_3/S FILL
XNOR3X1_1 NOR3X1_1/A INVX1_3/Y NOR3X1_1/C INVX1_3/gnd NOR3X1_1/Y DFFSR_79/S NOR3X1
XAND2X2_39 NOR2X1_70/A NOR2X1_70/B XOR2X1_4/gnd AND2X2_39/Y DFFSR_91/S AND2X2
XFILL_49_DFFSR_223 INVX1_39/gnd DFFSR_34/S FILL
XFILL_26_0_0 INVX1_3/gnd DFFSR_23/S FILL
XFILL_25_DFFSR_122 BUFX2_79/A DFFSR_7/S FILL
XFILL_38_DFFSR_37 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_39_DFFSR_226 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_1_INVX1_169 INVX1_39/gnd DFFSR_34/S FILL
XFILL_27_DFFSR_77 BUFX2_98/A DFFSR_32/S FILL
XFILL_4_AND2X2_36 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_15_DFFSR_125 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_7_NAND3X1_158 AND2X2_38/B DFFSR_59/S FILL
XFILL_29_DFFSR_229 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_5_AOI21X1_4 BUFX2_98/A DFFSR_32/S FILL
XFILL_24_2_1 AND2X2_38/B DFFSR_59/S FILL
XFILL_0_NAND2X1_139 INVX1_1/gnd DFFSR_97/S FILL
XDFFSR_34 DFFSR_34/Q AOI21X1_3/B DFFSR_1/R DFFSR_34/S DFFSR_34/D DFFSR_34/gnd DFFSR_34/S
+ DFFSR
XFILL_19_DFFSR_232 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_6_1_0 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_11_DFFSR_27 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_22_4_2 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_4_3_1 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_1_DFFSR_122 BUFX2_79/A DFFSR_7/S FILL
XFILL_42_DFFSR_153 INVX1_67/gnd DFFSR_201/S FILL
XFILL_51_1 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_46_DFFSR_44 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_35_DFFSR_84 BUFX2_99/A DFFSR_7/S FILL
XFILL_5_DFFSR_229 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_32_DFFSR_156 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_2_5_2 INVX1_67/gnd DFFSR_201/S FILL
XFILL_46_DFFSR_260 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_22_DFFSR_159 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_2_DFFSR_41 BUFX2_98/A DFFSR_6/S FILL
XFILL_36_DFFSR_263 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_19_DFFSR_34 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_7_NAND3X1_3 BUFX2_99/A DFFSR_92/S FILL
XFILL_12_DFFSR_162 BUFX2_99/A DFFSR_92/S FILL
XFILL_6_BUFX2_69 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_26_DFFSR_266 INVX1_67/gnd DFFSR_201/S FILL
XFILL_8_OAI21X1_110 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_16_DFFSR_269 INVX1_67/gnd DFFSR_201/S FILL
XFILL_6_NAND3X1_188 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_20_CLKBUF1_24 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_19_DFFSR_7 BUFX2_79/A DFFSR_7/S FILL
XFILL_12_XOR2X1_4 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_19_CLKBUF1_27 INVX1_1/gnd DFFSR_97/S FILL
XFILL_8_DFFSR_156 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_43_DFFSR_91 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_18_CLKBUF1_30 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_49_DFFSR_187 DFFSR_1/gnd DFFSR_81/S FILL
XNAND3X1_224 INVX1_169/Y AOI21X1_40/A AOI21X1_40/B INVX1_39/gnd AOI21X1_41/B DFFSR_54/S
+ NAND3X1
XFILL_17_CLKBUF1_33 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_1_INVX1_133 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_39_DFFSR_190 INVX1_39/gnd DFFSR_34/S FILL
XFILL_27_DFFSR_41 BUFX2_98/A DFFSR_6/S FILL
XFILL_16_DFFSR_81 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_2_DFFSR_266 INVX1_67/gnd DFFSR_201/S FILL
XFILL_7_NAND3X1_122 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_29_DFFSR_193 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_16_CLKBUF1_36 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_11_DFFPOSX1_26 AND2X2_38/B DFFSR_23/S FILL
XFILL_3_BUFX2_8 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_19_DFFSR_196 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_15_CLKBUF1_39 INVX1_1/gnd DFFSR_53/S FILL
XFILL_0_NAND2X1_103 AND2X2_38/B DFFSR_23/S FILL
XNOR2X1_78 XOR2X1_9/A XOR2X1_9/B NOR3X1_6/gnd NOR2X1_78/Y DFFSR_91/S NOR2X1
XFILL_14_CLKBUF1_42 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_51_DFFSR_98 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_13_CLKBUF1_45 BUFX2_79/A DFFSR_7/S FILL
XFILL_4_NOR2X1_75 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_40_DFFSR_3 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_12_CLKBUF1_48 INVX1_3/gnd DFFSR_79/S FILL
XFILL_21_DFFPOSX1_15 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_42_DFFSR_117 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_35_DFFSR_48 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_24_DFFSR_88 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_7_DFFSR_95 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_5_DFFSR_193 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_32_DFFSR_120 INVX1_3/gnd DFFSR_23/S FILL
XFILL_46_DFFSR_224 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_5_NAND3X1_218 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_22_DFFSR_123 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_1_DFFPOSX1_37 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_36_DFFSR_227 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_1_AND2X2_37 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_12_DFFSR_126 BUFX2_99/A DFFSR_7/S FILL
XFILL_6_BUFX2_33 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_26_DFFSR_230 INVX1_67/gnd DFFSR_201/S FILL
XFILL_2_AOI21X1_5 INVX1_3/gnd DFFSR_23/S FILL
XFILL_16_DFFSR_233 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_6_NAND3X1_152 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_43_DFFSR_55 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_32_DFFSR_95 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_8_DFFSR_120 INVX1_3/gnd DFFSR_23/S FILL
XFILL_49_DFFSR_151 XOR2X1_1/gnd DFFSR_151/S FILL
XNAND3X1_188 INVX1_157/A OAI21X1_59/C OAI21X1_52/Y BUFX2_7/gnd AOI21X1_26/B DFFSR_151/S
+ NAND3X1
XFILL_39_DFFSR_154 BUFX2_99/A DFFSR_7/S FILL
XFILL_16_DFFSR_45 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_2_DFFSR_230 INVX1_67/gnd DFFSR_201/S FILL
XFILL_3_BUFX2_80 BUFX2_79/A DFFSR_6/S FILL
XFILL_29_DFFSR_157 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_43_DFFSR_261 BUFX2_77/gnd DFFSR_98/S FILL
XNAND3X1_7 NAND3X1_7/A NAND3X1_7/B AOI22X1_1/Y OR2X2_6/gnd NOR2X1_8/B DFFSR_92/S NAND3X1
XFILL_19_DFFSR_160 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_20_DFFPOSX1_45 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_33_DFFSR_264 DFFSR_4/gnd DFFSR_98/S FILL
XNOR2X1_42 NOR2X1_42/A NOR2X1_42/B BUFX2_8/gnd NOR2X1_42/Y DFFSR_81/S NOR2X1
XFILL_4_NAND3X1_4 BUFX2_79/A DFFSR_7/S FILL
XFILL_23_DFFSR_267 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_4_NAND3X1_248 INVX1_3/gnd DFFSR_79/S FILL
XFILL_4_NOR2X1_39 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_13_DFFSR_270 INVX1_39/gnd DFFSR_54/S FILL
XFILL_12_CLKBUF1_12 AND2X2_38/B DFFSR_23/S FILL
XFILL_7_OAI21X1_104 INVX1_67/gnd DFFSR_201/S FILL
XFILL_35_DFFSR_12 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_24_DFFSR_52 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_7_DFFSR_59 AND2X2_38/B DFFSR_59/S FILL
XFILL_11_CLKBUF1_15 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_5_DFFSR_157 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_13_DFFSR_92 BUFX2_99/A DFFSR_92/S FILL
XFILL_23_5_0 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_46_DFFSR_188 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_10_CLKBUF1_18 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_5_NAND3X1_182 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_9_DFFSR_264 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_36_DFFSR_191 INVX1_67/gnd DFFSR_175/S FILL
XFILL_9_CLKBUF1_21 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_26_DFFSR_194 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_7_DFFSR_6 BUFX2_79/A DFFSR_6/S FILL
XFILL_16_DFFSR_197 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_8_CLKBUF1_24 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_3_6_0 INVX1_67/gnd DFFSR_175/S FILL
XFILL_6_NAND3X1_116 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_7_CLKBUF1_27 INVX1_1/gnd DFFSR_97/S FILL
XFILL_10_DFFPOSX1_20 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_43_DFFSR_19 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_4_INVX1_53 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_21_DFFSR_99 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_32_DFFSR_59 AND2X2_38/B DFFSR_59/S FILL
XFILL_6_CLKBUF1_30 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_1_NOR2X1_76 INVX1_3/gnd DFFSR_79/S FILL
XFILL_49_DFFSR_115 INVX1_1/gnd DFFSR_97/S FILL
XFILL_5_CLKBUF1_33 XOR2X1_4/gnd DFFSR_91/S FILL
XNAND3X1_152 INVX1_143/A NAND3X1_152/B NAND3X1_152/C DFFSR_34/gnd AOI21X1_9/B DFFSR_1/S
+ NAND3X1
XFILL_39_DFFSR_118 OR2X2_3/gnd DFFSR_60/S FILL
XCLKBUF1_30 BUFX2_2/Y BUFX2_77/gnd DFFSR_5/CLK DFFSR_5/S CLKBUF1
XFILL_5_OR2X2_6 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_4_CLKBUF1_36 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_2_DFFSR_194 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_3_BUFX2_44 INVX1_3/gnd DFFSR_79/S FILL
XFILL_29_DFFSR_121 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_43_DFFSR_225 INVX1_67/gnd DFFSR_175/S FILL
XFILL_3_CLKBUF1_39 INVX1_1/gnd DFFSR_53/S FILL
XFILL_8_AND2X2_35 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_19_DFFSR_124 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_2_CLKBUF1_42 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_33_DFFSR_228 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_9_AOI21X1_3 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_23_DFFSR_231 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_1_CLKBUF1_45 BUFX2_79/A DFFSR_7/S FILL
XFILL_4_NAND3X1_212 INVX1_39/gnd DFFSR_54/S FILL
XFILL_40_DFFSR_66 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_13_DFFSR_234 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_0_DFFPOSX1_31 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_0_CLKBUF1_48 INVX1_3/gnd DFFSR_79/S FILL
XFILL_16_3 INVX1_39/gnd DFFSR_34/S FILL
XFILL_33_0_0 INVX1_1/gnd DFFSR_53/S FILL
XFILL_24_DFFSR_16 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_7_DFFSR_23 AND2X2_38/B DFFSR_23/S FILL
XFILL_13_DFFSR_56 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_5_DFFSR_121 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_0_BUFX2_91 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_46_DFFSR_152 INVX1_1/gnd DFFSR_53/S FILL
XFILL_5_NAND3X1_146 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_31_2_1 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_9_DFFSR_228 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_36_DFFSR_155 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_6_NOR2X1_4 INVX1_1/gnd DFFSR_53/S FILL
XFILL_50_DFFSR_259 BUFX2_79/A DFFSR_6/S FILL
XFILL_26_DFFSR_158 INVX1_3/gnd DFFSR_23/S FILL
XFILL_40_DFFSR_262 BUFX2_98/A DFFSR_32/S FILL
XFILL_2_INVX1_205 BUFX2_99/A DFFSR_92/S FILL
XFILL_29_4_2 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_48_DFFSR_73 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_16_DFFSR_161 INVX1_67/gnd DFFSR_175/S FILL
XFILL_30_DFFSR_265 INVX1_67/gnd DFFSR_175/S FILL
XFILL_1_NAND3X1_5 BUFX2_99/A DFFSR_7/S FILL
XFILL_20_DFFSR_268 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_4_DFFSR_70 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_4_INVX1_17 AND2X2_38/B DFFSR_59/S FILL
XFILL_19_DFFPOSX1_39 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_21_DFFSR_63 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_32_DFFSR_23 AND2X2_38/B DFFSR_23/S FILL
XFILL_1_NOR2X1_40 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_10_DFFSR_271 BUFX2_8/gnd DFFSR_81/S FILL
XNAND3X1_116 NAND2X1_50/Y NAND3X1_113/Y AND2X2_25/Y DFFSR_46/gnd NOR2X1_55/A DFFSR_54/S
+ NAND3X1
XFILL_9_5_2 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_3_NAND3X1_242 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_2_DFFSR_158 INVX1_3/gnd DFFSR_23/S FILL
XFILL_43_DFFSR_189 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_6_DFFSR_265 INVX1_67/gnd DFFSR_175/S FILL
XFILL_33_DFFSR_192 INVX1_1/gnd DFFSR_97/S FILL
XFILL_4_NAND3X1_176 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_23_DFFSR_195 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_29_DFFSR_70 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_40_DFFSR_30 BUFX2_98/A DFFSR_32/S FILL
XFILL_1_INVX1_64 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_13_DFFSR_198 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_0_CLKBUF1_12 AND2X2_38/B DFFSR_23/S FILL
XFILL_9_DFFPOSX1_50 INVX1_1/gnd DFFSR_53/S FILL
XFILL_13_DFFSR_20 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_0_BUFX2_55 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_46_DFFSR_116 INVX1_3/gnd DFFSR_23/S FILL
XFILL_5_NAND3X1_110 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_9_DFFSR_192 INVX1_1/gnd DFFSR_97/S FILL
XFILL_36_DFFSR_119 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_4_NOR3X1_1 INVX1_3/gnd DFFSR_79/S FILL
XFILL_50_DFFSR_223 INVX1_39/gnd DFFSR_34/S FILL
XFILL_18_DFFSR_4 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_26_DFFSR_122 BUFX2_79/A DFFSR_7/S FILL
XFILL_40_DFFSR_226 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_2_INVX1_169 INVX1_39/gnd DFFSR_34/S FILL
XFILL_48_DFFSR_37 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_37_DFFSR_77 BUFX2_98/A DFFSR_32/S FILL
XFILL_5_AND2X2_36 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_16_DFFSR_125 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_30_DFFSR_229 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_6_AOI21X1_4 BUFX2_98/A DFFSR_32/S FILL
XFILL_20_DFFSR_232 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_4_DFFSR_34 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_21_DFFSR_27 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_10_DFFSR_67 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_2_BUFX2_5 AND2X2_38/B DFFSR_59/S FILL
XFILL_10_DFFSR_235 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_3_NAND3X1_206 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_2_DFFSR_122 BUFX2_79/A DFFSR_7/S FILL
XFILL_43_DFFSR_153 INVX1_67/gnd DFFSR_201/S FILL
XFILL_45_DFFSR_84 BUFX2_99/A DFFSR_7/S FILL
XFILL_6_DFFSR_229 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_33_DFFSR_156 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_47_DFFSR_260 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_4_NAND3X1_140 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_23_DFFSR_159 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_1_INVX1_28 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_37_DFFSR_263 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_1_DFFSR_81 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_29_DFFSR_34 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_18_DFFSR_74 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_8_NAND3X1_3 BUFX2_99/A DFFSR_92/S FILL
XFILL_13_DFFSR_162 BUFX2_99/A DFFSR_92/S FILL
XFILL_27_DFFSR_266 INVX1_67/gnd DFFSR_201/S FILL
XFILL_23_DFFPOSX1_3 INVX1_39/gnd DFFSR_34/S FILL
XFILL_9_DFFPOSX1_14 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_6_NAND2X1_176 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_17_DFFSR_269 INVX1_67/gnd DFFSR_201/S FILL
XFILL_22_DFFPOSX1_6 AND2X2_38/B DFFSR_23/S FILL
XFILL_0_BUFX2_19 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_21_DFFPOSX1_9 INVX1_67/gnd DFFSR_201/S FILL
XFILL_9_DFFSR_156 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_18_DFFPOSX1_33 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_50_DFFSR_187 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_2_INVX1_133 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_40_DFFSR_190 INVX1_39/gnd DFFSR_34/S FILL
XFILL_9_DFFSR_88 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_37_DFFSR_41 BUFX2_98/A DFFSR_6/S FILL
XFILL_26_DFFSR_81 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_2_NAND3X1_236 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_3_DFFSR_266 INVX1_67/gnd DFFSR_201/S FILL
XFILL_30_DFFSR_193 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_20_DFFSR_196 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_10_DFFSR_31 BUFX2_79/A DFFSR_6/S FILL
XFILL_10_DFFSR_199 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_30_5_0 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_5_NOR2X1_75 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_3_NAND3X1_170 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_18_NOR3X1_5 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_8_DFFPOSX1_44 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_43_DFFSR_117 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_45_DFFSR_48 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_6_DFFSR_193 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_34_DFFSR_88 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_33_DFFSR_120 INVX1_3/gnd DFFSR_23/S FILL
XFILL_47_DFFSR_224 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_23_DFFSR_123 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_4_NAND3X1_104 AND2X2_38/B DFFSR_23/S FILL
XFILL_37_DFFSR_227 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_1_DFFSR_45 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_18_DFFSR_38 BUFX2_98/A DFFSR_6/S FILL
XFILL_2_AND2X2_37 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_13_DFFSR_126 BUFX2_99/A DFFSR_7/S FILL
XFILL_5_BUFX2_73 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_27_DFFSR_230 INVX1_67/gnd DFFSR_201/S FILL
XFILL_6_NAND2X1_140 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_3_AOI21X1_5 INVX1_3/gnd DFFSR_23/S FILL
XFILL_17_DFFSR_233 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_6_DFFSR_3 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_11_XOR2X1_8 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_42_DFFSR_95 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_9_DFFSR_120 INVX1_3/gnd DFFSR_23/S FILL
XNAND2X1_176 XOR2X1_13/Y XOR2X1_14/Y XOR2X1_4/gnd AOI21X1_68/C DFFSR_97/S NAND2X1
XFILL_50_DFFSR_151 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_8_AOI21X1_68 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_3_AND2X2_4 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_40_DFFSR_154 BUFX2_99/A DFFSR_7/S FILL
XFILL_15_DFFSR_85 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_26_DFFSR_45 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_9_DFFSR_52 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_7_AOI21X1_71 BUFX2_99/A DFFSR_92/S FILL
XFILL_2_NAND3X1_200 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_3_DFFSR_230 INVX1_67/gnd DFFSR_201/S FILL
XFILL_30_DFFSR_157 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_44_DFFSR_261 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_20_DFFSR_160 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_4_OR2X2_3 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_34_DFFSR_264 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_40_0_0 BUFX2_98/A DFFSR_6/S FILL
XFILL_5_NAND3X1_4 BUFX2_79/A DFFSR_7/S FILL
XFILL_10_DFFSR_163 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_24_DFFSR_267 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_5_NOR2X1_39 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_3_NAND3X1_134 INVX1_39/gnd DFFSR_54/S FILL
XFILL_30_DFFSR_7 BUFX2_79/A DFFSR_7/S FILL
XFILL_38_2_1 BUFX2_79/A DFFSR_7/S FILL
XFILL_14_DFFSR_270 INVX1_39/gnd DFFSR_54/S FILL
XFILL_5_NAND2X1_170 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_45_DFFSR_12 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_34_DFFSR_52 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_6_DFFSR_99 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_6_DFFSR_157 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_23_DFFSR_92 BUFX2_99/A DFFSR_92/S FILL
XFILL_36_4_2 BUFX2_99/A DFFSR_92/S FILL
XFILL_47_DFFSR_188 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_11_DFFPOSX1_3 INVX1_39/gnd DFFSR_34/S FILL
XFILL_37_DFFSR_191 INVX1_67/gnd DFFSR_175/S FILL
XBUFX2_77 BUFX2_77/A BUFX2_77/gnd dout[6] DFFSR_5/S BUFX2
XFILL_5_BUFX2_37 INVX1_1/gnd DFFSR_97/S FILL
XFILL_10_DFFPOSX1_6 AND2X2_38/B DFFSR_23/S FILL
XFILL_0_DFFSR_267 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_27_DFFSR_194 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_17_DFFPOSX1_27 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_6_NAND2X1_104 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_17_DFFSR_197 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_1_NAND3X1_230 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_51_DFFSR_3 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_9_DFFPOSX1_9 INVX1_67/gnd DFFSR_201/S FILL
XFILL_31_DFFSR_99 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_3_INVX1_93 INVX1_3/gnd DFFSR_23/S FILL
XFILL_42_DFFSR_59 AND2X2_38/B DFFSR_59/S FILL
XNAND2X1_140 NAND2X1_143/A INVX1_208/Y BUFX2_7/gnd AOI21X1_46/A DFFSR_151/S NAND2X1
XFILL_2_NOR2X1_76 INVX1_3/gnd DFFSR_79/S FILL
XFILL_50_DFFSR_115 INVX1_1/gnd DFFSR_97/S FILL
XFILL_27_DFFPOSX1_16 INVX1_67/gnd DFFSR_175/S FILL
XFILL_8_AOI21X1_32 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_9_DFFSR_16 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_40_DFFSR_118 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_15_DFFSR_49 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_7_AOI21X1_35 INVX1_39/gnd DFFSR_54/S FILL
XFILL_3_DFFSR_194 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_2_NAND3X1_164 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_30_DFFSR_121 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_2_BUFX2_84 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_6_AOI21X1_38 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_44_DFFSR_225 INVX1_67/gnd DFFSR_175/S FILL
XFILL_20_DFFSR_124 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_7_DFFPOSX1_38 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_5_AOI21X1_41 INVX1_39/gnd DFFSR_34/S FILL
XFILL_34_DFFSR_228 XOR2X1_1/gnd DFFSR_208/S FILL
XAOI21X1_38 AOI21X1_38/A AOI21X1_38/B XOR2X1_8/B DFFSR_28/gnd AOI21X1_38/Y DFFSR_8/S
+ AOI21X1
XFILL_10_DFFSR_127 BUFX2_99/A DFFSR_92/S FILL
XFILL_4_AOI21X1_44 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_24_DFFSR_231 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_50_DFFSR_66 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_0_AOI21X1_6 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_3_AOI21X1_47 INVX1_67/gnd DFFSR_175/S FILL
XFILL_14_DFFSR_234 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_2_AOI21X1_50 INVX1_67/gnd DFFSR_175/S FILL
XFILL_34_DFFSR_16 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_6_DFFSR_63 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_5_NAND2X1_134 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_23_DFFSR_56 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_1_AOI21X1_53 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_12_DFFSR_96 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_6_DFFSR_121 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_47_DFFSR_152 INVX1_1/gnd DFFSR_53/S FILL
XFILL_0_AOI21X1_56 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_37_DFFSR_155 OR2X2_1/gnd DFFSR_59/S FILL
XBUFX2_41 INVX1_59/Y BUFX2_77/gnd DFFSR_35/R DFFSR_5/S BUFX2
XFILL_0_DFFSR_231 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_27_DFFSR_158 INVX1_3/gnd DFFSR_23/S FILL
XFILL_3_OAI21X1_116 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_41_DFFSR_262 BUFX2_98/A DFFSR_32/S FILL
XFILL_3_INVX1_205 BUFX2_99/A DFFSR_92/S FILL
XFILL_26_DFFPOSX1_46 INVX1_39/gnd DFFSR_34/S FILL
XFILL_17_DFFSR_161 INVX1_67/gnd DFFSR_175/S FILL
XFILL_31_DFFSR_265 INVX1_67/gnd DFFSR_175/S FILL
XFILL_8_OAI21X1_80 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_17_DFFSR_1 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_1_NAND3X1_194 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_2_NAND3X1_5 BUFX2_99/A DFFSR_7/S FILL
XFILL_7_OAI21X1_83 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_21_DFFSR_268 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_31_DFFSR_63 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_3_INVX1_57 BUFX2_98/A DFFSR_32/S FILL
XFILL_42_DFFSR_23 AND2X2_38/B DFFSR_23/S FILL
XNAND2X1_104 INVX1_133/A OR2X2_6/gnd OR2X2_6/gnd XOR2X1_5/A DFFSR_53/S NAND2X1
XFILL_2_NOR2X1_40 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_6_OAI21X1_86 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_11_DFFSR_271 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_12_0_1 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_5_OAI21X1_89 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_1_BUFX2_2 OR2X2_4/gnd DFFSR_32/S FILL
XOAI21X1_86 DFFSR_98/S INVX1_182/Y OAI21X1_86/C BUFX2_77/gnd DFFSR_258/D DFFSR_5/S
+ OAI21X1
XFILL_15_DFFSR_13 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_2_NAND3X1_128 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_3_DFFSR_158 INVX1_3/gnd DFFSR_23/S FILL
XFILL_4_OAI21X1_92 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_2_BUFX2_48 AND2X2_38/B DFFSR_59/S FILL
XFILL_44_DFFSR_189 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_3_OAI21X1_95 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_10_2_2 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_7_DFFSR_265 INVX1_67/gnd DFFSR_175/S FILL
XFILL_4_NAND2X1_164 INVX1_67/gnd DFFSR_175/S FILL
XFILL_34_DFFSR_192 INVX1_1/gnd DFFSR_97/S FILL
XFILL_2_OAI21X1_98 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_24_DFFSR_195 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_50_DFFSR_30 BUFX2_98/A DFFSR_32/S FILL
XFILL_39_DFFSR_70 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_3_AOI21X1_11 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_3_4 INVX1_67/gnd DFFSR_201/S FILL
XFILL_14_DFFSR_198 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_16_DFFPOSX1_21 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_2_AOI21X1_14 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_6_DFFSR_27 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_1_AOI21X1_17 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_12_DFFSR_60 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_23_DFFSR_20 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_0_NAND3X1_224 INVX1_39/gnd DFFSR_54/S FILL
XFILL_47_DFFSR_116 INVX1_3/gnd DFFSR_23/S FILL
XFILL_0_AOI21X1_20 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_37_DFFSR_119 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_5_NOR2X1_8 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_51_DFFSR_223 INVX1_39/gnd DFFSR_34/S FILL
XFILL_0_DFFSR_195 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_27_DFFSR_122 BUFX2_79/A DFFSR_7/S FILL
XFILL_26_DFFPOSX1_10 INVX1_67/gnd DFFSR_201/S FILL
XFILL_41_DFFSR_226 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_3_INVX1_169 INVX1_39/gnd DFFSR_34/S FILL
XFILL_47_DFFSR_77 BUFX2_98/A DFFSR_32/S FILL
XFILL_6_AND2X2_36 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_17_DFFSR_125 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_37_5_0 BUFX2_99/A DFFSR_7/S FILL
XFILL_31_DFFSR_229 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_8_OAI21X1_44 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_1_NAND3X1_158 AND2X2_38/B DFFSR_59/S FILL
XFILL_7_AOI21X1_4 BUFX2_98/A DFFSR_32/S FILL
XFILL_6_NAND2X1_65 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_7_OAI21X1_47 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_21_DFFSR_232 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_31_DFFSR_27 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_3_DFFSR_74 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_3_INVX1_21 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_20_DFFSR_67 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_6_DFFPOSX1_32 INVX1_67/gnd DFFSR_201/S FILL
XFILL_6_OAI21X1_50 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_5_NAND2X1_68 AND2X2_38/B DFFSR_23/S FILL
XFILL_11_DFFSR_235 OR2X2_2/gnd DFFSR_216/S FILL
XNAND2X1_65 AOI21X1_7/B AOI21X1_7/A XOR2X1_1/gnd NAND2X1_65/Y DFFSR_151/S NAND2X1
XFILL_4_NAND2X1_71 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_5_OAI21X1_53 XOR2X1_1/gnd DFFSR_151/S FILL
XOAI21X1_50 INVX1_132/Y INVX1_161/Y NOR2X1_70/A XOR2X1_4/gnd AOI21X1_30/B DFFSR_97/S
+ OAI21X1
XFILL_3_DFFSR_122 BUFX2_79/A DFFSR_7/S FILL
XFILL_2_BUFX2_12 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_3_NAND2X1_74 AND2X2_38/B DFFSR_59/S FILL
XFILL_4_OAI21X1_56 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_7_XOR2X1_4 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_44_DFFSR_153 INVX1_67/gnd DFFSR_201/S FILL
XFILL_2_NAND2X1_77 AND2X2_38/B DFFSR_23/S FILL
XFILL_3_OAI21X1_59 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_7_DFFSR_229 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_4_NAND2X1_128 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_34_DFFSR_156 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_2_OAI21X1_62 INVX1_3/gnd DFFSR_79/S FILL
XFILL_1_NAND2X1_80 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_48_DFFSR_260 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_11_AOI22X1_28 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_24_DFFSR_159 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_0_INVX1_68 INVX1_67/gnd DFFSR_201/S FILL
XFILL_1_OAI21X1_65 INVX1_1/gnd DFFSR_53/S FILL
XFILL_38_DFFSR_263 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_0_NAND2X1_83 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_28_DFFSR_74 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_0_INVX1_206 INVX1_1/gnd DFFSR_53/S FILL
XFILL_39_DFFSR_34 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_14_DFFSR_162 BUFX2_99/A DFFSR_92/S FILL
XFILL_28_DFFSR_266 INVX1_67/gnd DFFSR_201/S FILL
XFILL_0_OAI21X1_68 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_2_OAI21X1_110 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_18_DFFSR_269 INVX1_67/gnd DFFSR_201/S FILL
XFILL_25_DFFPOSX1_40 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_12_DFFSR_24 BUFX2_98/A DFFSR_6/S FILL
XFILL_0_NAND3X1_188 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_3_NOR3X1_5 BUFX2_7/gnd DFFSR_216/S FILL
XDFFSR_4 DFFSR_4/Q CLKBUF1_4/Y DFFSR_8/R DFFSR_4/S DFFSR_4/D DFFSR_4/gnd DFFSR_4/S
+ DFFSR
XDFFSR_269 INVX1_194/A CLKBUF1_47/Y DFFSR_266/R DFFSR_201/S DFFSR_269/D INVX1_67/gnd
+ DFFSR_201/S DFFSR
XFILL_47_0_0 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_0_DFFSR_159 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_3_INVX1_133 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_41_DFFSR_190 INVX1_39/gnd DFFSR_34/S FILL
XFILL_47_DFFSR_41 BUFX2_98/A DFFSR_6/S FILL
XFILL_36_DFFSR_81 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_4_DFFSR_266 INVX1_67/gnd DFFSR_201/S FILL
XFILL_31_DFFSR_193 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_1_NAND3X1_122 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_45_2_1 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_21_DFFSR_196 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_6_NAND2X1_29 INVX1_3/gnd DFFSR_23/S FILL
XFILL_7_OAI21X1_11 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_3_DFFSR_38 BUFX2_98/A DFFSR_6/S FILL
XFILL_20_DFFSR_31 BUFX2_79/A DFFSR_6/S FILL
XFILL_3_NAND2X1_158 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_5_NAND2X1_32 INVX1_3/gnd DFFSR_79/S FILL
XFILL_6_OAI21X1_14 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_11_DFFSR_199 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_43_4_2 OR2X2_4/gnd DFFSR_3/S FILL
XNAND2X1_29 NOR2X1_31/Y AND2X2_15/Y INVX1_3/gnd OAI22X1_41/D DFFSR_23/S NAND2X1
XFILL_4_NAND2X1_35 INVX1_67/gnd DFFSR_201/S FILL
XFILL_5_OAI21X1_17 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_6_NOR2X1_75 BUFX2_8/gnd DFFSR_51/S FILL
XOAI21X1_14 INVX1_103/Y OAI21X1_9/B NAND2X1_47/Y DFFSR_62/gnd NOR2X1_51/B DFFSR_208/S
+ OAI21X1
XFILL_4_OAI21X1_20 AND2X2_38/B DFFSR_23/S FILL
XFILL_3_NAND2X1_38 BUFX2_8/gnd DFFSR_81/S FILL
XDFFPOSX1_32 NAND2X1_163/B CLKBUF1_44/Y AOI21X1_58/Y INVX1_67/gnd DFFSR_201/S DFFPOSX1
XFILL_44_DFFSR_117 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_13_XOR2X1_1 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_15_DFFPOSX1_15 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_3_OAI21X1_23 INVX1_67/gnd DFFSR_201/S FILL
XFILL_2_NAND2X1_41 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_29_DFFSR_4 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_44_DFFSR_88 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_7_DFFSR_193 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_34_DFFSR_120 INVX1_3/gnd DFFSR_23/S FILL
XFILL_9_NAND3X1_97 AND2X2_38/B DFFSR_59/S FILL
XFILL_2_OAI21X1_26 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_1_NAND2X1_44 INVX1_39/gnd DFFSR_34/S FILL
XFILL_48_DFFSR_224 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_24_DFFSR_123 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_0_NAND2X1_47 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_1_OAI21X1_29 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_38_DFFSR_227 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_0_INVX1_32 OR2X2_6/gnd DFFSR_53/S FILL
XAOI21X1_8 AOI21X1_8/A AOI21X1_8/B NOR2X1_65/Y DFFSR_1/gnd AOI21X1_8/Y DFFSR_1/S AOI21X1
XFILL_0_INVX1_170 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_0_DFFSR_85 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_17_DFFSR_78 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_28_DFFSR_38 BUFX2_98/A DFFSR_6/S FILL
XFILL_3_AND2X2_37 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_14_DFFSR_126 BUFX2_99/A DFFSR_7/S FILL
XFILL_28_DFFSR_230 INVX1_67/gnd DFFSR_201/S FILL
XFILL_0_OAI21X1_32 AND2X2_38/B DFFSR_59/S FILL
XFILL_4_AOI21X1_5 INVX1_3/gnd DFFSR_23/S FILL
XFILL_11_3_0 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_18_DFFSR_233 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_0_NAND3X1_152 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_5_DFFPOSX1_26 AND2X2_38/B DFFSR_23/S FILL
XDFFSR_233 DFFSR_241/D CLKBUF1_2/Y BUFX2_62/Y DFFSR_175/S DFFSR_225/Q OR2X2_2/gnd
+ DFFSR_175/S DFFSR
XFILL_0_DFFSR_123 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_41_DFFSR_154 BUFX2_99/A DFFSR_7/S FILL
XFILL_36_DFFSR_45 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_8_DFFSR_92 BUFX2_99/A DFFSR_92/S FILL
XFILL_25_DFFSR_85 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_4_DFFSR_230 INVX1_67/gnd DFFSR_201/S FILL
XFILL_5_AOI22X1_10 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_31_DFFSR_157 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_45_DFFSR_261 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_4_AOI22X1_13 AND2X2_38/B DFFSR_23/S FILL
XFILL_21_DFFSR_160 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_35_DFFSR_264 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_14_DFFPOSX1_45 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_3_AOI22X1_16 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_3_NAND2X1_122 INVX1_67/gnd DFFSR_175/S FILL
XFILL_6_NAND3X1_4 BUFX2_79/A DFFSR_7/S FILL
XFILL_11_DFFSR_163 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_2_AOI22X1_19 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_25_DFFSR_267 XOR2X1_1/gnd DFFSR_208/S FILL
XINVX1_6 INVX1_6/A BUFX2_8/gnd INVX1_6/Y DFFSR_81/S INVX1
XFILL_6_NOR2X1_39 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_15_DFFSR_270 INVX1_39/gnd DFFSR_54/S FILL
XFILL_11_OAI22X1_40 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_1_AOI22X1_22 INVX1_3/gnd DFFSR_79/S FILL
XFILL_0_AOI22X1_25 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_10_OAI22X1_43 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_1_OAI21X1_104 INVX1_67/gnd DFFSR_201/S FILL
XFILL_7_DFFSR_157 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_44_DFFSR_52 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_33_DFFSR_92 BUFX2_99/A DFFSR_92/S FILL
XFILL_24_DFFPOSX1_34 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_48_DFFSR_188 DFFSR_46/gnd DFFSR_54/S FILL
XAND2X2_1 INVX1_3/Y NOR3X1_1/A XOR2X1_4/gnd AND2X2_1/Y DFFSR_97/S AND2X2
XFILL_8_NAND3X1_64 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_0_NAND2X1_11 BUFX2_98/A DFFSR_6/S FILL
XFILL_9_OAI22X1_46 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_38_DFFSR_191 INVX1_67/gnd DFFSR_175/S FILL
XFILL_8_NAND3X1_237 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_0_INVX1_134 INVX1_3/gnd DFFSR_79/S FILL
XFILL_17_DFFSR_42 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_0_DFFSR_49 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_7_NAND3X1_67 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_4_BUFX2_77 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_8_OAI22X1_49 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_1_DFFSR_267 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_28_DFFSR_194 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_6_NAND3X1_70 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_7_OAI22X1_52 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_18_DFFSR_197 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_19_0_1 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_5_NAND3X1_73 INVX1_1/gnd DFFSR_97/S FILL
XFILL_0_NAND3X1_116 DFFSR_46/gnd DFFSR_54/S FILL
XNAND3X1_70 DFFSR_201/D BUFX2_28/Y NOR2X1_31/Y BUFX2_7/gnd NAND3X1_71/B DFFSR_151/S
+ NAND3X1
XFILL_4_NAND3X1_76 INVX1_1/gnd DFFSR_53/S FILL
XFILL_41_DFFSR_99 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_9_NAND3X1_171 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_3_NOR2X1_76 INVX1_3/gnd DFFSR_79/S FILL
XFILL_17_2_2 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_3_NAND3X1_79 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_2_NAND2X1_152 INVX1_1/gnd DFFSR_97/S FILL
XDFFSR_197 DFFSR_205/D CLKBUF1_40/Y BUFX2_63/Y DFFSR_97/S DFFSR_141/Q XOR2X1_4/gnd
+ DFFSR_97/S DFFSR
XFILL_41_DFFSR_118 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_2_AND2X2_8 BUFX2_99/A DFFSR_7/S FILL
XFILL_2_NAND3X1_82 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_8_DFFSR_56 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_25_DFFSR_49 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_14_DFFSR_89 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_4_DFFSR_194 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_31_DFFSR_121 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_1_NAND3X1_85 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_45_DFFSR_225 INVX1_67/gnd DFFSR_175/S FILL
XFILL_21_DFFSR_124 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_0_NAND3X1_88 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_35_DFFSR_228 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_0_AND2X2_38 AND2X2_38/B DFFSR_59/S FILL
XFILL_11_DFFSR_127 BUFX2_99/A DFFSR_92/S FILL
XFILL_25_DFFSR_231 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_1_AOI21X1_6 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_15_DFFSR_234 OR2X2_3/gnd DFFSR_4/S FILL
XINVX1_90 INVX1_90/A NOR3X1_6/gnd INVX1_90/Y DFFSR_79/S INVX1
XFILL_44_DFFSR_16 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_33_DFFSR_56 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_22_DFFSR_96 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_7_DFFSR_121 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_44_5_0 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_48_DFFSR_152 INVX1_1/gnd DFFSR_53/S FILL
XFILL_8_NAND3X1_28 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_9_OAI22X1_10 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_0_DFFSR_13 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_8_NAND3X1_201 INVX1_1/gnd DFFSR_53/S FILL
XFILL_38_DFFSR_155 OR2X2_1/gnd DFFSR_59/S FILL
XINVX1_208 DFFSR_54/S INVX1_39/gnd INVX1_208/Y DFFSR_34/S INVX1
XFILL_4_BUFX2_41 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_7_NAND3X1_31 BUFX2_79/A DFFSR_6/S FILL
XFILL_8_OAI22X1_13 INVX1_1/gnd DFFSR_53/S FILL
XFILL_1_DFFSR_231 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_28_DFFSR_158 INVX1_3/gnd DFFSR_23/S FILL
XFILL_4_DFFPOSX1_20 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_42_DFFSR_262 BUFX2_98/A DFFSR_32/S FILL
XFILL_1_NAND2X1_182 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_6_NAND3X1_34 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_4_INVX1_205 BUFX2_99/A DFFSR_92/S FILL
XFILL_7_OAI22X1_16 AND2X2_38/B DFFSR_59/S FILL
XFILL_18_DFFSR_161 INVX1_67/gnd DFFSR_175/S FILL
XFILL_32_DFFSR_265 INVX1_67/gnd DFFSR_175/S FILL
XFILL_6_OAI22X1_19 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_5_NAND3X1_37 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_41_DFFSR_7 BUFX2_79/A DFFSR_7/S FILL
XFILL_3_NAND3X1_5 BUFX2_99/A DFFSR_7/S FILL
XNAND3X1_34 DFFSR_5/Q NOR2X1_4/Y BUFX2_15/Y DFFSR_8/gnd AND2X2_10/B DFFSR_60/S NAND3X1
XFILL_22_DFFSR_268 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_5_OAI22X1_22 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_41_DFFSR_63 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_4_NAND3X1_40 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_2_INVX1_97 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_3_NOR2X1_40 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_13_DFFPOSX1_39 BUFX2_7/gnd DFFSR_151/S FILL
XOAI22X1_19 INVX1_45/Y OAI22X1_7/B INVX1_46/Y OAI22X1_7/D OR2X2_3/gnd NOR2X1_24/B
+ DFFSR_60/S OAI22X1
XFILL_12_DFFSR_271 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_3_NAND3X1_43 BUFX2_99/A DFFSR_7/S FILL
XFILL_4_OAI22X1_25 INVX1_39/gnd DFFSR_54/S FILL
XDFFSR_161 DFFSR_161/Q CLKBUF1_2/Y BUFX2_67/Y DFFSR_175/S INVX1_66/A INVX1_67/gnd
+ DFFSR_175/S DFFSR
XFILL_2_NAND2X1_116 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_2_NAND3X1_46 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_3_OAI22X1_28 INVX1_3/gnd DFFSR_23/S FILL
XFILL_8_DFFSR_20 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_25_DFFSR_13 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_14_DFFSR_53 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_4_DFFSR_158 INVX1_3/gnd DFFSR_23/S FILL
XFILL_1_NAND3X1_49 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_1_BUFX2_88 INVX1_3/gnd DFFSR_23/S FILL
XFILL_2_OAI22X1_31 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_45_DFFSR_189 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_8_DFFSR_265 INVX1_67/gnd DFFSR_175/S FILL
XFILL_0_NAND3X1_52 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_1_OAI22X1_34 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_35_DFFSR_192 INVX1_1/gnd DFFSR_97/S FILL
XFILL_23_DFFPOSX1_28 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_0_OAI22X1_37 INVX1_3/gnd DFFSR_23/S FILL
XFILL_25_DFFSR_195 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_49_DFFSR_70 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_7_1 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_15_DFFSR_198 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_7_NAND3X1_231 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_3_DFFPOSX1_50 INVX1_1/gnd DFFSR_53/S FILL
XFILL_54_0_0 DFFSR_5/gnd DFFSR_5/S FILL
XINVX1_54 INVX1_54/A DFFSR_4/gnd INVX1_54/Y DFFSR_4/S INVX1
XFILL_22_DFFSR_60 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_33_DFFSR_20 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_5_DFFSR_67 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_0_NOR2X1_77 INVX1_39/gnd DFFSR_34/S FILL
XFILL_48_DFFSR_116 INVX1_3/gnd DFFSR_23/S FILL
XFILL_52_2_1 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_38_DFFSR_119 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_8_NAND3X1_165 INVX1_39/gnd DFFSR_34/S FILL
XINVX1_172 INVX1_172/A DFFSR_28/gnd XOR2X1_8/B DFFSR_8/S INVX1
XFILL_1_DFFSR_195 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_28_DFFSR_122 BUFX2_79/A DFFSR_7/S FILL
XFILL_1_NAND2X1_146 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_42_DFFSR_226 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_4_INVX1_169 INVX1_39/gnd DFFSR_34/S FILL
XFILL_18_DFFSR_125 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_7_AND2X2_36 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_50_4_2 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_32_DFFSR_229 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_8_AOI21X1_4 BUFX2_98/A DFFSR_32/S FILL
XFILL_22_DFFSR_232 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_41_DFFSR_27 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_2_INVX1_61 INVX1_39/gnd DFFSR_54/S FILL
XFILL_30_DFFSR_67 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_12_DFFSR_235 OR2X2_2/gnd DFFSR_216/S FILL
XDFFSR_125 BUFX2_86/A DFFSR_93/CLK DFFSR_5/R DFFSR_5/S INVX1_37/A DFFSR_5/gnd DFFSR_5/S
+ DFFSR
XFILL_2_NAND3X1_10 BUFX2_79/A DFFSR_6/S FILL
XFILL_14_DFFSR_17 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_4_DFFSR_122 BUFX2_79/A DFFSR_7/S FILL
XFILL_1_BUFX2_52 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_1_NAND3X1_13 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_45_DFFSR_153 INVX1_67/gnd DFFSR_201/S FILL
XFILL_0_NAND3X1_16 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_8_DFFSR_229 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_35_DFFSR_156 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_18_3_0 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_49_DFFSR_260 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_28_DFFSR_1 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_25_DFFSR_159 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_39_DFFSR_263 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_38_DFFSR_74 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_1_INVX1_206 INVX1_1/gnd DFFSR_53/S FILL
XFILL_49_DFFSR_34 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_15_DFFSR_162 BUFX2_99/A DFFSR_92/S FILL
XFILL_16_5_1 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_7_NAND3X1_195 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_29_DFFSR_266 INVX1_67/gnd DFFSR_201/S FILL
XFILL_0_NAND3X1_6 BUFX2_99/A DFFSR_92/S FILL
XFILL_3_DFFPOSX1_14 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_19_DFFSR_269 INVX1_67/gnd DFFSR_201/S FILL
XFILL_0_NAND2X1_176 XOR2X1_4/gnd DFFSR_97/S FILL
XDFFSR_71 DFFSR_79/D DFFSR_79/CLK DFFSR_7/R DFFSR_91/S DFFSR_71/D XOR2X1_4/gnd DFFSR_91/S
+ DFFSR
XINVX1_18 DFFSR_51/D OR2X2_1/gnd INVX1_18/Y DFFSR_59/S INVX1
XFILL_11_DFFSR_64 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_22_DFFSR_24 BUFX2_98/A DFFSR_6/S FILL
XFILL_5_DFFSR_31 BUFX2_79/A DFFSR_6/S FILL
XFILL_0_NOR2X1_41 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_8_NAND3X1_129 DFFSR_62/gnd DFFSR_62/S FILL
XINVX1_136 INVX1_136/A OR2X2_2/gnd OR2X2_2/B DFFSR_216/S INVX1
XFILL_12_DFFPOSX1_33 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_1_DFFSR_159 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_1_NAND2X1_110 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_4_INVX1_133 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_42_DFFSR_190 INVX1_39/gnd DFFSR_34/S FILL
XFILL_46_DFFSR_81 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_5_DFFSR_266 INVX1_67/gnd DFFSR_201/S FILL
XFILL_32_DFFSR_193 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_22_DFFSR_196 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_2_INVX1_25 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_2_DFFSR_78 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_30_DFFSR_31 BUFX2_79/A DFFSR_6/S FILL
XFILL_19_DFFSR_71 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_12_DFFSR_199 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_22_DFFPOSX1_22 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_6_NAND3X1_225 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_1_BUFX2_16 BUFX2_98/A DFFSR_32/S FILL
XFILL_6_XOR2X1_8 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_45_DFFSR_117 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_2_DFFPOSX1_44 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_8_DFFSR_193 OR2X2_2/gnd DFFSR_175/S FILL
XNOR3X1_2 OR2X2_1/A BUFX2_9/Y NOR3X1_2/C INVX1_1/gnd NOR3X1_2/Y DFFSR_53/S NOR3X1
XFILL_35_DFFSR_120 INVX1_3/gnd DFFSR_23/S FILL
XFILL_49_DFFSR_224 BUFX2_7/gnd DFFSR_151/S FILL
XAND2X2_40 AND2X2_40/A INVX1_180/Y OR2X2_4/gnd AND2X2_40/Y DFFSR_32/S AND2X2
XFILL_26_0_1 INVX1_3/gnd DFFSR_23/S FILL
XFILL_25_DFFSR_123 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_39_DFFSR_227 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_1_INVX1_170 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_27_DFFSR_78 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_38_DFFSR_38 BUFX2_98/A DFFSR_6/S FILL
XFILL_4_AND2X2_37 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_15_DFFSR_126 BUFX2_99/A DFFSR_7/S FILL
XFILL_7_NAND3X1_159 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_29_DFFSR_230 INVX1_67/gnd DFFSR_201/S FILL
XFILL_5_AOI21X1_5 INVX1_3/gnd DFFSR_23/S FILL
XFILL_24_2_2 AND2X2_38/B DFFSR_59/S FILL
XFILL_19_DFFSR_233 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_0_NAND2X1_140 BUFX2_7/gnd DFFSR_151/S FILL
XDFFSR_35 DFFSR_43/D DFFSR_57/CLK DFFSR_35/R DFFSR_3/S INVX1_21/A DFFSR_28/gnd DFFSR_3/S
+ DFFSR
XFILL_11_DFFSR_28 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_6_1_1 BUFX2_7/gnd DFFSR_216/S FILL
XINVX1_100 DFFSR_214/D OR2X2_2/gnd INVX1_100/Y DFFSR_175/S INVX1
XFILL_4_3_2 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_1_DFFSR_123 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_42_DFFSR_154 BUFX2_99/A DFFSR_7/S FILL
XFILL_46_DFFSR_45 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_51_2 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_35_DFFSR_85 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_5_DFFSR_230 INVX1_67/gnd DFFSR_201/S FILL
XFILL_32_DFFSR_157 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_46_DFFSR_261 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_22_DFFSR_160 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_36_DFFSR_264 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_2_DFFSR_42 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_19_DFFSR_35 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_7_NAND3X1_4 BUFX2_79/A DFFSR_7/S FILL
XFILL_6_BUFX2_70 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_12_DFFSR_163 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_26_DFFSR_267 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_8_OAI21X1_111 AND2X2_38/B DFFSR_59/S FILL
XFILL_51_5_0 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_16_DFFSR_270 INVX1_39/gnd DFFSR_54/S FILL
XFILL_20_CLKBUF1_25 INVX1_67/gnd DFFSR_201/S FILL
XFILL_6_NAND3X1_189 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_12_XOR2X1_5 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_19_DFFSR_8 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_19_CLKBUF1_28 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_43_DFFSR_92 BUFX2_99/A DFFSR_92/S FILL
XFILL_8_DFFSR_157 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_18_CLKBUF1_31 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_49_DFFSR_188 DFFSR_46/gnd DFFSR_54/S FILL
XNAND3X1_225 OAI21X1_77/Y INVX1_177/Y NAND2X1_107/Y DFFSR_4/gnd NAND3X1_227/A DFFSR_4/S
+ NAND3X1
XFILL_4_AND2X2_1 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_17_CLKBUF1_34 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_39_DFFSR_191 INVX1_67/gnd DFFSR_175/S FILL
XFILL_27_DFFSR_42 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_1_INVX1_134 INVX1_3/gnd DFFSR_79/S FILL
XFILL_16_DFFSR_82 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_7_NAND3X1_123 BUFX2_99/A DFFSR_7/S FILL
XFILL_2_DFFSR_267 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_29_DFFSR_194 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_16_CLKBUF1_37 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_3_BUFX2_9 AND2X2_38/B DFFSR_59/S FILL
XFILL_11_DFFPOSX1_27 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_0_NAND2X1_104 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_15_CLKBUF1_40 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_19_DFFSR_197 XOR2X1_4/gnd DFFSR_97/S FILL
XNOR2X1_79 BUFX2_39/Y NOR2X1_79/B DFFSR_46/gnd NOR2X1_79/Y DFFSR_54/S NOR2X1
XFILL_14_CLKBUF1_43 AND2X2_38/B DFFSR_23/S FILL
XFILL_13_CLKBUF1_46 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_40_DFFSR_4 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_4_NOR2X1_76 INVX1_3/gnd DFFSR_79/S FILL
XFILL_12_CLKBUF1_49 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_21_DFFPOSX1_16 INVX1_67/gnd DFFSR_175/S FILL
XFILL_42_DFFSR_118 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_7_DFFSR_96 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_35_DFFSR_49 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_24_DFFSR_89 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_5_DFFSR_194 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_32_DFFSR_121 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_46_DFFSR_225 INVX1_67/gnd DFFSR_175/S FILL
XFILL_5_NAND3X1_219 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_22_DFFSR_124 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_36_DFFSR_228 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_1_DFFPOSX1_38 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_1_AND2X2_38 AND2X2_38/B DFFSR_59/S FILL
XFILL_12_DFFSR_127 BUFX2_99/A DFFSR_92/S FILL
XFILL_6_BUFX2_34 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_26_DFFSR_231 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_2_AOI21X1_6 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_16_DFFSR_234 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_6_NAND3X1_153 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_43_DFFSR_56 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_32_DFFSR_96 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_4_INVX1_90 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_8_DFFSR_121 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_49_DFFSR_152 INVX1_1/gnd DFFSR_53/S FILL
XNAND3X1_189 INVX1_157/Y OAI21X1_53/Y OAI21X1_54/Y BUFX2_7/gnd AOI21X1_26/A DFFSR_151/S
+ NAND3X1
XFILL_39_DFFSR_155 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_16_DFFSR_46 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_2_DFFSR_231 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_3_BUFX2_81 BUFX2_79/A DFFSR_7/S FILL
XFILL_29_DFFSR_158 INVX1_3/gnd DFFSR_23/S FILL
XFILL_43_DFFSR_262 BUFX2_98/A DFFSR_32/S FILL
XNAND3X1_8 NOR2X1_3/Y NOR2X1_6/Y NOR2X1_8/Y XOR2X1_4/gnd NAND3X1_8/Y DFFSR_97/S NAND3X1
XFILL_20_DFFPOSX1_46 INVX1_39/gnd DFFSR_34/S FILL
XFILL_19_DFFSR_161 INVX1_67/gnd DFFSR_175/S FILL
XFILL_33_DFFSR_265 INVX1_67/gnd DFFSR_175/S FILL
XFILL_4_NAND3X1_5 BUFX2_99/A DFFSR_7/S FILL
XNOR2X1_43 NOR2X1_43/A NOR2X1_43/B DFFSR_34/gnd NOR2X1_43/Y DFFSR_34/S NOR2X1
XFILL_4_NAND3X1_249 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_23_DFFSR_268 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_51_DFFSR_63 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_13_CLKBUF1_10 INVX1_67/gnd DFFSR_201/S FILL
XFILL_4_NOR2X1_40 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_13_DFFSR_271 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_25_3_0 AND2X2_38/B DFFSR_23/S FILL
XFILL_12_CLKBUF1_13 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_7_OAI21X1_105 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_7_DFFSR_60 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_13_DFFSR_93 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_11_CLKBUF1_16 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_35_DFFSR_13 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_24_DFFSR_53 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_5_DFFSR_158 INVX1_3/gnd DFFSR_23/S FILL
XFILL_5_NAND3X1_183 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_23_5_1 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_46_DFFSR_189 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_10_CLKBUF1_19 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_9_DFFSR_265 INVX1_67/gnd DFFSR_175/S FILL
XFILL_36_DFFSR_192 INVX1_1/gnd DFFSR_97/S FILL
XFILL_5_4_0 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_9_CLKBUF1_22 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_26_DFFSR_195 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_7_DFFSR_7 BUFX2_79/A DFFSR_7/S FILL
XFILL_8_CLKBUF1_25 INVX1_67/gnd DFFSR_201/S FILL
XFILL_16_DFFSR_198 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_3_6_1 INVX1_67/gnd DFFSR_175/S FILL
XFILL_6_NAND3X1_117 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_7_CLKBUF1_28 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_10_DFFPOSX1_21 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_32_DFFSR_60 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_4_INVX1_54 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_43_DFFSR_20 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_6_CLKBUF1_31 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_1_NOR2X1_77 INVX1_39/gnd DFFSR_34/S FILL
XFILL_49_DFFSR_116 INVX1_3/gnd DFFSR_23/S FILL
XFILL_5_CLKBUF1_34 BUFX2_72/gnd DFFSR_201/S FILL
XNAND3X1_153 AOI21X1_9/C AOI21X1_9/A AOI21X1_9/B XOR2X1_1/gnd NOR3X1_5/A DFFSR_151/S
+ NAND3X1
XFILL_39_DFFSR_119 OR2X2_4/gnd DFFSR_3/S FILL
XCLKBUF1_31 BUFX2_3/Y BUFX2_72/gnd CLKBUF1_31/Y DFFSR_201/S CLKBUF1
XFILL_16_DFFSR_10 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_4_CLKBUF1_37 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_2_DFFSR_195 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_3_BUFX2_45 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_29_DFFSR_122 BUFX2_79/A DFFSR_7/S FILL
XFILL_43_DFFSR_226 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_3_CLKBUF1_40 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_20_DFFPOSX1_10 INVX1_67/gnd DFFSR_201/S FILL
XFILL_8_AND2X2_36 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_19_DFFSR_125 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_2_CLKBUF1_43 AND2X2_38/B DFFSR_23/S FILL
XFILL_33_DFFSR_229 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_9_AOI21X1_4 BUFX2_98/A DFFSR_32/S FILL
XFILL_1_CLKBUF1_46 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_4_NAND3X1_213 INVX1_39/gnd DFFSR_54/S FILL
XFILL_23_DFFSR_232 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_51_DFFSR_27 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_40_DFFSR_67 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_0_DFFPOSX1_32 INVX1_67/gnd DFFSR_201/S FILL
XFILL_13_DFFSR_235 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_0_CLKBUF1_49 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_16_4 INVX1_39/gnd DFFSR_34/S FILL
XFILL_33_0_1 INVX1_1/gnd DFFSR_53/S FILL
XFILL_7_DFFSR_24 BUFX2_98/A DFFSR_6/S FILL
XFILL_24_DFFSR_17 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_13_DFFSR_57 BUFX2_79/A DFFSR_6/S FILL
XFILL_5_DFFSR_122 BUFX2_79/A DFFSR_7/S FILL
XFILL_0_BUFX2_92 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_46_DFFSR_153 INVX1_67/gnd DFFSR_201/S FILL
XFILL_5_NAND3X1_147 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_31_2_2 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_9_DFFSR_229 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_36_DFFSR_156 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_50_DFFSR_260 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_6_NOR2X1_5 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_26_DFFSR_159 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_40_DFFSR_263 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_48_DFFSR_74 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_2_INVX1_206 INVX1_1/gnd DFFSR_53/S FILL
XFILL_16_DFFSR_162 BUFX2_99/A DFFSR_92/S FILL
XFILL_30_DFFSR_266 INVX1_67/gnd DFFSR_201/S FILL
XFILL_1_NAND3X1_6 BUFX2_99/A DFFSR_92/S FILL
XFILL_20_DFFSR_269 INVX1_67/gnd DFFSR_201/S FILL
XFILL_32_DFFSR_24 BUFX2_98/A DFFSR_6/S FILL
XFILL_4_DFFSR_71 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_21_DFFSR_64 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_19_DFFPOSX1_40 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_1_NOR2X1_41 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_10_DFFSR_272 INVX1_3/gnd DFFSR_23/S FILL
XNAND3X1_117 DFFSR_143/Q BUFX2_31/Y BUFX2_24/Y DFFSR_62/gnd NAND3X1_117/Y DFFSR_208/S
+ NAND3X1
XFILL_3_NAND3X1_243 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_2_DFFSR_159 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_8_XOR2X1_1 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_43_DFFSR_190 INVX1_39/gnd DFFSR_34/S FILL
XFILL_6_DFFSR_266 INVX1_67/gnd DFFSR_201/S FILL
XFILL_33_DFFSR_193 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_1_CLKBUF1_10 INVX1_67/gnd DFFSR_201/S FILL
XFILL_23_DFFSR_196 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_4_NAND3X1_177 AND2X2_38/B DFFSR_59/S FILL
XFILL_1_INVX1_65 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_40_DFFSR_31 BUFX2_79/A DFFSR_6/S FILL
XFILL_29_DFFSR_71 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_0_CLKBUF1_13 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_13_DFFSR_199 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_13_DFFSR_21 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_0_BUFX2_56 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_5_NAND3X1_111 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_46_DFFSR_117 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_9_DFFSR_193 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_36_DFFSR_120 INVX1_3/gnd DFFSR_23/S FILL
XFILL_4_NOR3X1_2 INVX1_1/gnd DFFSR_53/S FILL
XFILL_50_DFFSR_224 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_18_DFFSR_5 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_26_DFFSR_123 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_40_DFFSR_227 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_2_INVX1_170 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_37_DFFSR_78 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_48_DFFSR_38 BUFX2_98/A DFFSR_6/S FILL
XFILL_5_AND2X2_37 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_16_DFFSR_126 BUFX2_99/A DFFSR_7/S FILL
XFILL_30_DFFSR_230 INVX1_67/gnd DFFSR_201/S FILL
XFILL_6_AOI21X1_5 INVX1_3/gnd DFFSR_23/S FILL
XFILL_20_DFFSR_233 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_4_DFFSR_35 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_21_DFFSR_28 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_10_DFFSR_68 BUFX2_98/A DFFSR_6/S FILL
XFILL_2_BUFX2_6 BUFX2_79/A DFFSR_6/S FILL
XFILL_10_DFFSR_236 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_3_NAND3X1_207 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_2_DFFSR_123 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_43_DFFSR_154 BUFX2_99/A DFFSR_7/S FILL
XFILL_39_DFFSR_1 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_45_DFFSR_85 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_6_DFFSR_230 INVX1_67/gnd DFFSR_201/S FILL
XFILL_33_DFFSR_157 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_47_DFFSR_261 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_23_DFFSR_160 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_4_NAND3X1_141 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_29_DFFSR_35 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_1_INVX1_29 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_37_DFFSR_264 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_1_DFFSR_82 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_18_DFFSR_75 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_8_NAND3X1_4 BUFX2_79/A DFFSR_7/S FILL
XFILL_24_DFFPOSX1_1 INVX1_39/gnd DFFSR_34/S FILL
XFILL_13_DFFSR_163 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_27_DFFSR_267 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_9_DFFPOSX1_15 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_23_DFFPOSX1_4 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_6_NAND2X1_177 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_17_DFFSR_270 INVX1_39/gnd DFFSR_54/S FILL
XFILL_22_DFFPOSX1_7 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_0_BUFX2_20 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_9_DFFSR_157 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_18_DFFPOSX1_34 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_50_DFFSR_188 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_40_DFFSR_191 INVX1_67/gnd DFFSR_175/S FILL
XFILL_37_DFFSR_42 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_2_INVX1_134 INVX1_3/gnd DFFSR_79/S FILL
XFILL_9_DFFSR_89 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_26_DFFSR_82 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_2_NAND3X1_237 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_3_DFFSR_267 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_30_DFFSR_194 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_32_3_0 INVX1_1/gnd DFFSR_97/S FILL
XFILL_20_DFFSR_197 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_10_DFFSR_32 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_10_DFFSR_200 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_30_5_1 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_5_NOR2X1_76 INVX1_3/gnd DFFSR_79/S FILL
XFILL_3_NAND3X1_171 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_18_NOR3X1_6 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_43_DFFSR_118 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_8_DFFPOSX1_45 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_45_DFFSR_49 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_34_DFFSR_89 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_6_DFFSR_194 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_33_DFFSR_121 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_47_DFFSR_225 INVX1_67/gnd DFFSR_175/S FILL
XFILL_23_DFFSR_124 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_4_NAND3X1_105 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_18_DFFSR_39 INVX1_3/gnd DFFSR_79/S FILL
XFILL_1_DFFSR_46 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_37_DFFSR_228 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_2_AND2X2_38 AND2X2_38/B DFFSR_59/S FILL
XFILL_5_BUFX2_74 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_13_DFFSR_127 BUFX2_99/A DFFSR_92/S FILL
XFILL_27_DFFSR_231 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_3_AOI21X1_6 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_6_NAND2X1_141 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_17_DFFSR_234 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_6_DFFSR_4 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_11_XOR2X1_9 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_42_DFFSR_96 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_9_DFFSR_121 OR2X2_6/gnd DFFSR_53/S FILL
XNAND2X1_177 XOR2X1_13/Y AOI21X1_67/A XOR2X1_4/gnd OAI21X1_116/C DFFSR_97/S NAND2X1
XFILL_50_DFFSR_152 INVX1_1/gnd DFFSR_53/S FILL
XFILL_8_AOI21X1_69 INVX1_1/gnd DFFSR_97/S FILL
XFILL_3_AND2X2_5 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_40_DFFSR_155 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_9_DFFSR_53 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_15_DFFSR_86 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_26_DFFSR_46 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_2_NAND3X1_201 INVX1_1/gnd DFFSR_53/S FILL
XFILL_3_DFFSR_231 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_30_DFFSR_158 INVX1_3/gnd DFFSR_23/S FILL
XFILL_44_DFFSR_262 BUFX2_98/A DFFSR_32/S FILL
XFILL_20_DFFSR_161 INVX1_67/gnd DFFSR_175/S FILL
XFILL_4_OR2X2_4 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_34_DFFSR_265 INVX1_67/gnd DFFSR_175/S FILL
XFILL_40_0_1 BUFX2_98/A DFFSR_6/S FILL
XFILL_5_NAND3X1_5 BUFX2_99/A DFFSR_7/S FILL
XFILL_10_DFFSR_164 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_24_DFFSR_268 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_5_NOR2X1_40 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_3_NAND3X1_135 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_30_DFFSR_8 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_14_DFFSR_271 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_38_2_2 BUFX2_79/A DFFSR_7/S FILL
XFILL_23_DFFSR_93 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_45_DFFSR_13 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_34_DFFSR_53 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_5_NAND2X1_171 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_6_DFFSR_158 INVX1_3/gnd DFFSR_23/S FILL
XFILL_12_DFFPOSX1_1 INVX1_39/gnd DFFSR_34/S FILL
XFILL_47_DFFSR_189 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_11_DFFPOSX1_4 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_1_DFFSR_10 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_37_DFFSR_192 INVX1_1/gnd DFFSR_97/S FILL
XFILL_10_DFFPOSX1_7 OR2X2_3/gnd DFFSR_4/S FILL
XBUFX2_78 BUFX2_78/A DFFSR_4/gnd dout[7] DFFSR_4/S BUFX2
XFILL_0_DFFSR_268 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_5_BUFX2_38 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_17_DFFPOSX1_28 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_27_DFFSR_195 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_6_NAND2X1_105 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_17_DFFSR_198 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_1_NAND3X1_231 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_3_INVX1_94 INVX1_67/gnd DFFSR_201/S FILL
XFILL_42_DFFSR_60 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_2_NOR2X1_77 INVX1_39/gnd DFFSR_34/S FILL
XNAND2X1_141 NAND2X1_144/A DFFSR_54/S DFFSR_46/gnd AOI21X1_46/B DFFSR_62/S NAND2X1
XFILL_50_DFFSR_116 INVX1_3/gnd DFFSR_23/S FILL
XFILL_8_AOI21X1_33 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_27_DFFPOSX1_17 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_40_DFFSR_119 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_9_DFFSR_17 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_7_AOI21X1_36 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_26_DFFSR_10 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_15_DFFSR_50 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_2_NAND3X1_165 INVX1_39/gnd DFFSR_34/S FILL
XFILL_3_DFFSR_195 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_2_BUFX2_85 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_30_DFFSR_122 BUFX2_79/A DFFSR_7/S FILL
XFILL_6_AOI21X1_39 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_44_DFFSR_226 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_7_DFFPOSX1_39 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_20_DFFSR_125 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_5_AOI21X1_42 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_34_DFFSR_229 OR2X2_1/gnd DFFSR_59/S FILL
XAOI21X1_39 AOI21X1_39/A AOI21X1_39/B INVX1_172/A DFFSR_8/gnd OAI21X1_82/A DFFSR_8/S
+ AOI21X1
XFILL_10_DFFSR_128 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_4_AOI21X1_45 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_24_DFFSR_232 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_0_AOI21X1_7 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_50_DFFSR_67 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_14_DFFSR_235 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_20_1 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_3_AOI21X1_48 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_2_AOI21X1_51 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_34_DFFSR_17 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_6_DFFSR_64 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_23_DFFSR_57 BUFX2_79/A DFFSR_6/S FILL
XFILL_5_NAND2X1_135 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_6_DFFSR_122 BUFX2_79/A DFFSR_7/S FILL
XFILL_12_DFFSR_97 INVX1_1/gnd DFFSR_97/S FILL
XFILL_1_AOI21X1_54 AND2X2_38/B DFFSR_59/S FILL
XFILL_47_DFFSR_153 INVX1_67/gnd DFFSR_201/S FILL
XFILL_0_AOI21X1_57 INVX1_67/gnd DFFSR_201/S FILL
XFILL_37_DFFSR_156 OR2X2_2/gnd DFFSR_175/S FILL
XBUFX2_42 INVX1_59/Y OR2X2_4/gnd DFFSR_3/R DFFSR_3/S BUFX2
XFILL_0_DFFSR_232 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_3_OAI21X1_117 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_27_DFFSR_159 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_9_OAI21X1_78 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_3_INVX1_206 INVX1_1/gnd DFFSR_53/S FILL
XFILL_26_DFFPOSX1_47 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_41_DFFSR_263 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_17_DFFSR_162 BUFX2_99/A DFFSR_92/S FILL
XFILL_8_OAI21X1_81 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_17_DFFSR_2 BUFX2_79/A DFFSR_7/S FILL
XFILL_31_DFFSR_266 INVX1_67/gnd DFFSR_201/S FILL
XFILL_1_NAND3X1_195 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_2_NAND3X1_6 BUFX2_99/A DFFSR_92/S FILL
XFILL_21_DFFSR_269 INVX1_67/gnd DFFSR_201/S FILL
XFILL_7_OAI21X1_84 BUFX2_98/A DFFSR_6/S FILL
XFILL_42_DFFSR_24 BUFX2_98/A DFFSR_6/S FILL
XFILL_3_INVX1_58 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_31_DFFSR_64 OR2X2_3/gnd DFFSR_60/S FILL
XNAND2X1_105 AND2X2_35/A OR2X2_6/gnd OR2X2_6/gnd XOR2X1_5/B DFFSR_53/S NAND2X1
XFILL_2_NOR2X1_41 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_6_OAI21X1_87 BUFX2_79/A DFFSR_7/S FILL
XFILL_11_DFFSR_272 INVX1_3/gnd DFFSR_23/S FILL
XFILL_5_OAI21X1_90 BUFX2_98/A DFFSR_32/S FILL
XFILL_12_0_2 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_1_BUFX2_3 BUFX2_8/gnd DFFSR_81/S FILL
XOAI21X1_87 DFFSR_7/S INVX1_183/Y OAI21X1_87/C BUFX2_79/A DFFSR_259/D DFFSR_7/S OAI21X1
XFILL_15_DFFSR_14 INVX1_1/gnd DFFSR_53/S FILL
XFILL_2_NAND3X1_129 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_4_OAI21X1_93 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_3_DFFSR_159 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_2_BUFX2_49 INVX1_1/gnd DFFSR_97/S FILL
XFILL_44_DFFSR_190 INVX1_39/gnd DFFSR_34/S FILL
XFILL_3_OAI21X1_96 AND2X2_38/B DFFSR_59/S FILL
XFILL_7_DFFSR_266 INVX1_67/gnd DFFSR_201/S FILL
XFILL_4_NAND2X1_165 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_34_DFFSR_193 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_2_OAI21X1_99 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_24_DFFSR_196 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_50_DFFSR_31 BUFX2_79/A DFFSR_6/S FILL
XFILL_39_DFFSR_71 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_3_AOI21X1_12 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_14_DFFSR_199 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_2_AOI21X1_15 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_16_DFFPOSX1_22 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_6_DFFSR_28 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_23_DFFSR_21 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_1_AOI21X1_18 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_12_DFFSR_61 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_0_DFFPOSX1_1 INVX1_39/gnd DFFSR_34/S FILL
XFILL_0_NAND3X1_225 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_47_DFFSR_117 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_0_AOI21X1_21 INVX1_39/gnd DFFSR_54/S FILL
XFILL_37_DFFSR_120 INVX1_3/gnd DFFSR_23/S FILL
XFILL_39_3_0 BUFX2_79/A DFFSR_6/S FILL
XFILL_5_NOR2X1_9 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_0_DFFSR_196 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_27_DFFSR_123 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_9_OAI21X1_42 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_26_DFFPOSX1_11 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_41_DFFSR_227 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_3_INVX1_170 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_47_DFFSR_78 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_6_AND2X2_37 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_17_DFFSR_126 BUFX2_99/A DFFSR_7/S FILL
XFILL_37_5_1 BUFX2_99/A DFFSR_7/S FILL
XFILL_8_OAI21X1_45 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_31_DFFSR_230 INVX1_67/gnd DFFSR_201/S FILL
XFILL_1_NAND3X1_159 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_7_AOI21X1_5 INVX1_3/gnd DFFSR_23/S FILL
XFILL_6_NAND2X1_66 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_21_DFFSR_233 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_7_OAI21X1_48 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_3_INVX1_22 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_31_DFFSR_28 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_20_DFFSR_68 BUFX2_98/A DFFSR_6/S FILL
XFILL_3_DFFSR_75 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_6_DFFPOSX1_33 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_5_NAND2X1_69 INVX1_3/gnd DFFSR_23/S FILL
XFILL_11_DFFSR_236 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_6_OAI21X1_51 DFFSR_62/gnd DFFSR_208/S FILL
XNAND2X1_66 INVX1_133/A INVX1_159/A BUFX2_8/gnd INVX1_143/A DFFSR_81/S NAND2X1
XFILL_4_NAND2X1_72 AND2X2_38/B DFFSR_59/S FILL
XFILL_5_OAI21X1_54 XOR2X1_1/gnd DFFSR_208/S FILL
XOAI21X1_51 OAI21X1_53/A OAI21X1_53/B OAI21X1_54/C DFFSR_62/gnd OAI21X1_59/C DFFSR_208/S
+ OAI21X1
XFILL_42_1 BUFX2_98/A DFFSR_32/S FILL
XFILL_3_DFFSR_123 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_3_NAND2X1_75 INVX1_3/gnd DFFSR_79/S FILL
XFILL_4_OAI21X1_57 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_2_BUFX2_13 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_44_DFFSR_154 BUFX2_99/A DFFSR_7/S FILL
XFILL_7_XOR2X1_5 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_10_AOI22X1_1 INVX1_1/gnd DFFSR_97/S FILL
XFILL_2_NAND2X1_78 AND2X2_38/B DFFSR_23/S FILL
XFILL_3_OAI21X1_60 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_7_DFFSR_230 INVX1_67/gnd DFFSR_201/S FILL
XFILL_4_NAND2X1_129 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_34_DFFSR_157 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_2_OAI21X1_63 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_1_NAND2X1_81 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_48_DFFSR_261 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_11_AOI22X1_29 INVX1_1/gnd DFFSR_53/S FILL
XFILL_24_DFFSR_160 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_1_OAI21X1_66 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_0_NAND2X1_84 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_39_DFFSR_35 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_38_DFFSR_264 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_0_INVX1_69 INVX1_3/gnd DFFSR_23/S FILL
XFILL_0_INVX1_207 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_28_DFFSR_75 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_14_DFFSR_163 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_0_OAI21X1_69 INVX1_3/gnd DFFSR_23/S FILL
XFILL_28_DFFSR_267 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_2_OAI21X1_111 AND2X2_38/B DFFSR_59/S FILL
XFILL_25_DFFPOSX1_41 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_18_DFFSR_270 INVX1_39/gnd DFFSR_54/S FILL
XFILL_12_DFFSR_25 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_0_NAND3X1_189 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_9_NAND3X1_244 DFFSR_28/gnd DFFSR_8/S FILL
XDFFSR_5 DFFSR_5/Q DFFSR_5/CLK DFFSR_5/R DFFSR_5/S DFFSR_5/D DFFSR_5/gnd DFFSR_5/S
+ DFFSR
XFILL_5_DFFSR_1 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_3_NOR3X1_6 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_51_DFFSR_188 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_0_DFFSR_160 XOR2X1_4/gnd DFFSR_97/S FILL
XDFFSR_270 INVX1_195/A CLKBUF1_44/Y DFFSR_266/R DFFSR_54/S DFFSR_270/D INVX1_39/gnd
+ DFFSR_54/S DFFSR
XFILL_47_0_1 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_41_DFFSR_191 INVX1_67/gnd DFFSR_175/S FILL
XFILL_3_INVX1_134 INVX1_3/gnd DFFSR_79/S FILL
XFILL_36_DFFSR_82 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_47_DFFSR_42 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_4_DFFSR_267 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_1_NAND3X1_123 BUFX2_99/A DFFSR_7/S FILL
XFILL_31_DFFSR_194 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_45_2_2 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_6_NAND2X1_30 AND2X2_38/B DFFSR_23/S FILL
XFILL_21_DFFSR_197 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_7_OAI21X1_12 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_3_DFFSR_39 INVX1_3/gnd DFFSR_79/S FILL
XFILL_20_DFFSR_32 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_3_NAND2X1_159 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_5_NAND2X1_33 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_6_OAI21X1_15 INVX1_3/gnd DFFSR_79/S FILL
XFILL_11_DFFSR_200 DFFSR_62/gnd DFFSR_62/S FILL
XNAND2X1_30 NOR2X1_30/Y NOR2X1_31/Y AND2X2_38/B OAI22X1_41/B DFFSR_23/S NAND2X1
XFILL_3_OR2X2_1 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_4_NAND2X1_36 INVX1_3/gnd DFFSR_79/S FILL
XFILL_5_OAI21X1_18 INVX1_39/gnd DFFSR_34/S FILL
XFILL_6_NOR2X1_76 INVX1_3/gnd DFFSR_79/S FILL
XOAI21X1_15 INVX1_110/Y OAI21X1_9/B OAI21X1_15/C INVX1_3/gnd NOR2X1_54/B DFFSR_79/S
+ OAI21X1
XFILL_3_NAND2X1_39 BUFX2_98/A DFFSR_6/S FILL
XFILL_4_OAI21X1_21 AND2X2_38/B DFFSR_59/S FILL
XDFFPOSX1_33 NAND2X1_157/B CLKBUF1_45/Y AOI21X1_55/Y XOR2X1_4/gnd DFFSR_91/S DFFPOSX1
XFILL_13_XOR2X1_2 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_44_DFFSR_118 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_29_DFFSR_5 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_15_DFFPOSX1_16 INVX1_67/gnd DFFSR_175/S FILL
XFILL_44_DFFSR_89 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_3_OAI21X1_24 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_2_NAND2X1_42 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_7_DFFSR_194 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_34_DFFSR_121 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_48_DFFSR_225 INVX1_67/gnd DFFSR_175/S FILL
XFILL_2_OAI21X1_27 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_1_NAND2X1_45 INVX1_39/gnd DFFSR_34/S FILL
XFILL_13_1_0 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_24_DFFSR_124 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_0_NAND2X1_48 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_1_OAI21X1_30 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_0_INVX1_33 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_0_DFFSR_86 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_0_INVX1_171 BUFX2_98/A DFFSR_6/S FILL
XFILL_28_DFFSR_39 INVX1_3/gnd DFFSR_79/S FILL
XFILL_38_DFFSR_228 XOR2X1_1/gnd DFFSR_208/S FILL
XAOI21X1_9 AOI21X1_9/A AOI21X1_9/B AOI21X1_9/C XOR2X1_1/gnd INVX1_147/A DFFSR_151/S
+ AOI21X1
XFILL_17_DFFSR_79 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_3_AND2X2_38 AND2X2_38/B DFFSR_59/S FILL
XFILL_14_DFFSR_127 BUFX2_99/A DFFSR_92/S FILL
XFILL_0_OAI21X1_33 INVX1_3/gnd DFFSR_79/S FILL
XFILL_28_DFFSR_231 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_4_AOI21X1_6 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_11_3_1 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_18_DFFSR_234 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_0_NAND3X1_153 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_9_NAND3X1_208 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_50_DFFSR_1 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_51_DFFSR_152 INVX1_1/gnd DFFSR_53/S FILL
XFILL_5_DFFPOSX1_27 DFFSR_34/gnd DFFSR_1/S FILL
XDFFSR_234 DFFSR_242/D DFFSR_5/CLK BUFX2_65/Y DFFSR_4/S DFFSR_234/D OR2X2_3/gnd DFFSR_4/S
+ DFFSR
XFILL_0_DFFSR_124 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_41_DFFSR_155 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_8_DFFSR_93 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_25_DFFSR_86 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_36_DFFSR_46 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_5_AOI22X1_11 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_4_DFFSR_231 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_31_DFFSR_158 INVX1_3/gnd DFFSR_23/S FILL
XFILL_4_AOI22X1_14 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_45_DFFSR_262 BUFX2_98/A DFFSR_32/S FILL
XFILL_21_DFFSR_161 INVX1_67/gnd DFFSR_175/S FILL
XFILL_14_DFFPOSX1_46 INVX1_39/gnd DFFSR_34/S FILL
XFILL_35_DFFSR_265 INVX1_67/gnd DFFSR_175/S FILL
XFILL_6_NAND3X1_5 BUFX2_99/A DFFSR_7/S FILL
XFILL_3_AOI22X1_17 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_11_DFFSR_164 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_3_NAND2X1_123 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_25_DFFSR_268 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_2_AOI22X1_20 INVX1_39/gnd DFFSR_34/S FILL
XINVX1_7 INVX1_7/A OR2X2_4/gnd INVX1_7/Y DFFSR_32/S INVX1
XFILL_6_NOR2X1_40 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_15_DFFSR_271 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_1_AOI22X1_23 INVX1_39/gnd DFFSR_34/S FILL
XFILL_11_OAI22X1_41 INVX1_39/gnd DFFSR_54/S FILL
XFILL_10_OAI22X1_44 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_0_AOI22X1_26 INVX1_1/gnd DFFSR_97/S FILL
XFILL_44_DFFSR_53 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_1_OAI21X1_105 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_33_DFFSR_93 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_7_DFFSR_158 INVX1_3/gnd DFFSR_23/S FILL
XFILL_24_DFFPOSX1_35 INVX1_39/gnd DFFSR_54/S FILL
XFILL_9_NAND3X1_62 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_48_DFFSR_189 BUFX2_8/gnd DFFSR_51/S FILL
XAND2X2_2 INVX1_4/Y BUFX2_7/Y BUFX2_99/A AND2X2_2/Y DFFSR_7/S AND2X2
XFILL_9_OAI22X1_47 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_8_NAND3X1_65 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_0_NAND2X1_12 INVX1_3/gnd DFFSR_79/S FILL
XFILL_0_DFFSR_50 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_8_NAND3X1_238 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_38_DFFSR_192 INVX1_1/gnd DFFSR_97/S FILL
XFILL_0_INVX1_135 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_17_DFFSR_43 BUFX2_98/A DFFSR_6/S FILL
XFILL_7_NAND3X1_68 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_4_BUFX2_78 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_8_OAI22X1_50 INVX1_3/gnd DFFSR_23/S FILL
XFILL_1_DFFSR_268 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_28_DFFSR_195 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_6_NAND3X1_71 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_18_DFFSR_198 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_19_0_2 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_5_NAND3X1_74 INVX1_1/gnd DFFSR_97/S FILL
XFILL_0_NAND3X1_117 DFFSR_62/gnd DFFSR_208/S FILL
XNAND3X1_71 NAND3X1_71/A NAND3X1_71/B AOI22X1_9/Y BUFX2_7/gnd NOR2X1_37/B DFFSR_216/S
+ NAND3X1
XFILL_4_NAND3X1_77 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_9_NAND3X1_172 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_3_NOR2X1_77 INVX1_39/gnd DFFSR_34/S FILL
XDFFSR_198 DFFSR_206/D CLKBUF1_21/Y BUFX2_68/Y DFFSR_216/S DFFSR_198/D BUFX2_7/gnd
+ DFFSR_216/S DFFSR
XFILL_3_NAND3X1_80 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_2_NAND2X1_153 BUFX2_98/A DFFSR_32/S FILL
XFILL_41_DFFSR_119 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_2_AND2X2_9 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_2_NAND3X1_83 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_36_DFFSR_10 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_25_DFFSR_50 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_14_DFFSR_90 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_8_DFFSR_57 BUFX2_79/A DFFSR_6/S FILL
XFILL_10_XNOR2X1_1 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_4_DFFSR_195 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_31_DFFSR_122 BUFX2_79/A DFFSR_7/S FILL
XFILL_1_NAND3X1_86 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_45_DFFSR_226 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_21_DFFSR_125 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_0_NAND3X1_89 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_14_DFFPOSX1_10 INVX1_67/gnd DFFSR_201/S FILL
XFILL_35_DFFSR_229 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_0_AND2X2_39 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_11_DFFSR_128 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_25_DFFSR_232 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_1_AOI21X1_7 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_15_DFFSR_235 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_46_3_0 DFFSR_8/gnd DFFSR_8/S FILL
XINVX1_91 INVX1_91/A AND2X2_38/B INVX1_91/Y DFFSR_23/S INVX1
XFILL_44_DFFSR_17 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_33_DFFSR_57 BUFX2_79/A DFFSR_6/S FILL
XFILL_7_DFFSR_122 BUFX2_79/A DFFSR_7/S FILL
XFILL_22_DFFSR_97 INVX1_1/gnd DFFSR_97/S FILL
XFILL_48_DFFSR_153 INVX1_67/gnd DFFSR_201/S FILL
XFILL_44_5_1 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_8_NAND3X1_29 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_9_OAI22X1_11 BUFX2_99/A DFFSR_92/S FILL
XFILL_38_DFFSR_156 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_8_NAND3X1_202 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_0_DFFSR_14 INVX1_1/gnd DFFSR_53/S FILL
XINVX1_209 NOR3X1_6/A NOR3X1_6/gnd INVX1_209/Y DFFSR_91/S INVX1
XFILL_8_OAI22X1_14 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_7_NAND3X1_32 BUFX2_79/A DFFSR_7/S FILL
XFILL_1_DFFSR_232 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_4_BUFX2_42 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_4_DFFPOSX1_21 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_28_DFFSR_159 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_4_INVX1_206 INVX1_1/gnd DFFSR_53/S FILL
XFILL_42_DFFSR_263 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_6_NAND3X1_35 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_7_OAI22X1_17 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_18_DFFSR_162 BUFX2_99/A DFFSR_92/S FILL
XFILL_32_DFFSR_266 INVX1_67/gnd DFFSR_201/S FILL
XFILL_41_DFFSR_8 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_6_OAI22X1_20 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_5_NAND3X1_38 BUFX2_98/A DFFSR_32/S FILL
XFILL_3_NAND3X1_6 BUFX2_99/A DFFSR_92/S FILL
XFILL_22_DFFSR_269 INVX1_67/gnd DFFSR_201/S FILL
XNAND3X1_35 BUFX2_86/A AND2X2_3/Y BUFX2_20/Y DFFSR_8/gnd AND2X2_10/A DFFSR_8/S NAND3X1
XFILL_5_OAI22X1_23 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_4_NAND3X1_41 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_41_DFFSR_64 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_2_INVX1_98 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_3_NOR2X1_41 DFFSR_1/gnd DFFSR_81/S FILL
XOAI22X1_20 INVX1_47/Y OAI22X1_2/B INVX1_48/Y OAI22X1_2/D DFFSR_4/gnd NOR2X1_24/A
+ DFFSR_98/S OAI22X1
XFILL_13_DFFPOSX1_40 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_3_NAND3X1_44 BUFX2_99/A DFFSR_7/S FILL
XFILL_12_DFFSR_272 INVX1_3/gnd DFFSR_23/S FILL
XDFFSR_162 DFFSR_170/D CLKBUF1_3/Y BUFX2_63/Y DFFSR_92/S INVX1_73/A BUFX2_99/A DFFSR_92/S
+ DFFSR
XFILL_4_OAI22X1_26 INVX1_39/gnd DFFSR_54/S FILL
XFILL_2_NAND2X1_117 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_2_NAND3X1_47 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_8_DFFSR_21 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_3_OAI22X1_29 INVX1_3/gnd DFFSR_79/S FILL
XFILL_25_DFFSR_14 INVX1_1/gnd DFFSR_53/S FILL
XFILL_14_DFFSR_54 INVX1_39/gnd DFFSR_54/S FILL
XFILL_4_DFFSR_159 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_1_NAND3X1_50 BUFX2_98/A DFFSR_6/S FILL
XFILL_1_BUFX2_89 INVX1_1/gnd DFFSR_97/S FILL
XFILL_2_OAI22X1_32 INVX1_39/gnd DFFSR_54/S FILL
XFILL_45_DFFSR_190 INVX1_39/gnd DFFSR_34/S FILL
XFILL_10_6_0 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_8_DFFSR_266 INVX1_67/gnd DFFSR_201/S FILL
XFILL_0_NAND3X1_53 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_1_OAI22X1_35 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_35_DFFSR_193 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_23_DFFPOSX1_29 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_0_OAI22X1_38 AND2X2_38/B DFFSR_23/S FILL
XFILL_25_DFFSR_196 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_49_DFFSR_71 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_7_2 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_15_DFFSR_199 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_7_NAND3X1_232 DFFSR_4/gnd DFFSR_98/S FILL
XINVX1_55 DFFSR_80/Q DFFSR_4/gnd INVX1_55/Y DFFSR_98/S INVX1
XFILL_54_0_1 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_33_DFFSR_21 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_5_DFFSR_68 BUFX2_98/A DFFSR_6/S FILL
XFILL_22_DFFSR_61 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_0_NOR2X1_78 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_48_DFFSR_117 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_52_2_2 BUFX2_77/gnd DFFSR_98/S FILL
XINVX1_173 XOR2X1_6/Y DFFSR_4/gnd INVX1_173/Y DFFSR_98/S INVX1
XFILL_38_DFFSR_120 INVX1_3/gnd DFFSR_23/S FILL
XFILL_8_NAND3X1_166 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_1_DFFSR_196 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_28_DFFSR_123 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_1_NAND2X1_147 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_42_DFFSR_227 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_7_AND2X2_37 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_18_DFFSR_126 BUFX2_99/A DFFSR_7/S FILL
XFILL_32_DFFSR_230 INVX1_67/gnd DFFSR_201/S FILL
XFILL_8_AOI21X1_5 INVX1_3/gnd DFFSR_23/S FILL
XFILL_22_DFFSR_233 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_41_DFFSR_28 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_30_DFFSR_68 BUFX2_98/A DFFSR_6/S FILL
XFILL_2_INVX1_62 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_12_DFFSR_236 DFFSR_62/gnd DFFSR_62/S FILL
XDFFSR_126 BUFX2_87/A CLKBUF1_40/Y BUFX2_49/Y DFFSR_7/S INVX1_44/A BUFX2_99/A DFFSR_7/S
+ DFFSR
XFILL_2_NAND3X1_11 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_20_1_0 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_14_DFFSR_18 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_4_DFFSR_123 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_1_BUFX2_53 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_1_NAND3X1_14 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_45_DFFSR_154 BUFX2_99/A DFFSR_7/S FILL
XFILL_11_AOI22X1_1 INVX1_1/gnd DFFSR_97/S FILL
XFILL_8_DFFSR_230 INVX1_67/gnd DFFSR_201/S FILL
XFILL_0_NAND3X1_17 BUFX2_99/A DFFSR_7/S FILL
XFILL_18_3_1 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_35_DFFSR_157 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_49_DFFSR_261 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_28_DFFSR_2 BUFX2_79/A DFFSR_7/S FILL
XFILL_25_DFFSR_160 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_0_2_0 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_49_DFFSR_35 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_39_DFFSR_264 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_1_INVX1_207 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_38_DFFSR_75 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_15_DFFSR_163 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_16_5_2 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_7_NAND3X1_196 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_29_DFFSR_267 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_0_NAND3X1_7 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_3_DFFPOSX1_15 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_0_NAND2X1_177 XOR2X1_4/gnd DFFSR_97/S FILL
XINVX1_19 DFFSR_83/Q NOR3X1_6/gnd INVX1_19/Y DFFSR_91/S INVX1
XFILL_19_DFFSR_270 INVX1_39/gnd DFFSR_54/S FILL
XDFFSR_72 DFFSR_72/Q CLKBUF1_5/Y DFFSR_35/R DFFSR_60/S DFFSR_16/Q OR2X2_3/gnd DFFSR_60/S
+ DFFSR
XFILL_5_DFFSR_32 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_22_DFFSR_25 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_11_DFFSR_65 BUFX2_79/A DFFSR_7/S FILL
XFILL_0_NOR2X1_42 BUFX2_8/gnd DFFSR_81/S FILL
XINVX1_137 INVX1_137/A OR2X2_2/gnd XOR2X1_2/B DFFSR_175/S INVX1
XFILL_8_NAND3X1_130 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_1_DFFSR_160 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_12_DFFPOSX1_34 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_1_NAND2X1_111 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_42_DFFSR_191 INVX1_67/gnd DFFSR_175/S FILL
XFILL_4_INVX1_134 INVX1_3/gnd DFFSR_79/S FILL
XFILL_46_DFFSR_82 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_5_DFFSR_267 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_32_DFFSR_194 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_22_DFFSR_197 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_30_DFFSR_32 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_2_INVX1_26 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_2_DFFSR_79 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_19_DFFSR_72 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_12_DFFSR_200 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_22_DFFPOSX1_23 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_1_BUFX2_17 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_6_NAND3X1_226 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_45_DFFSR_118 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_6_XOR2X1_9 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_2_DFFPOSX1_45 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_8_DFFSR_194 DFFSR_1/gnd DFFSR_81/S FILL
XNOR3X1_3 NOR3X1_3/A NOR3X1_3/B NOR3X1_3/C BUFX2_7/gnd NOR3X1_3/Y DFFSR_216/S NOR3X1
XFILL_35_DFFSR_121 OR2X2_6/gnd DFFSR_53/S FILL
XAND2X2_41 XOR2X1_9/Y NOR2X1_77/A DFFSR_1/gnd OR2X2_5/A DFFSR_81/S AND2X2
XFILL_49_DFFSR_225 INVX1_67/gnd DFFSR_175/S FILL
XFILL_26_0_2 INVX1_3/gnd DFFSR_23/S FILL
XFILL_25_DFFSR_124 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_1_INVX1_171 BUFX2_98/A DFFSR_6/S FILL
XFILL_39_DFFSR_228 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_27_DFFSR_79 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_38_DFFSR_39 INVX1_3/gnd DFFSR_79/S FILL
XFILL_4_AND2X2_38 AND2X2_38/B DFFSR_59/S FILL
XFILL_15_DFFSR_127 BUFX2_99/A DFFSR_92/S FILL
XFILL_7_NAND3X1_160 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_29_DFFSR_231 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_5_AOI21X1_6 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_19_DFFSR_234 OR2X2_3/gnd DFFSR_4/S FILL
XDFFSR_36 DFFSR_44/D CLKBUF1_37/Y DFFSR_8/R DFFSR_98/S INVX1_28/A BUFX2_77/gnd DFFSR_98/S
+ DFFSR
XFILL_0_NAND2X1_141 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_11_DFFSR_29 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_6_1_2 BUFX2_7/gnd DFFSR_216/S FILL
XINVX1_101 INVX1_101/A OR2X2_1/gnd INVX1_101/Y DFFSR_51/S INVX1
XFILL_1_DFFSR_124 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_42_DFFSR_155 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_51_3 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_35_DFFSR_86 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_46_DFFSR_46 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_5_DFFSR_231 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_32_DFFSR_158 INVX1_3/gnd DFFSR_23/S FILL
XFILL_46_DFFSR_262 BUFX2_98/A DFFSR_32/S FILL
XFILL_22_DFFSR_161 INVX1_67/gnd DFFSR_175/S FILL
XFILL_53_3_0 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_36_DFFSR_265 INVX1_67/gnd DFFSR_175/S FILL
XFILL_19_DFFSR_36 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_2_DFFSR_43 BUFX2_98/A DFFSR_6/S FILL
XFILL_12_DFFSR_164 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_7_NAND3X1_5 BUFX2_99/A DFFSR_7/S FILL
XFILL_6_BUFX2_71 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_26_DFFSR_268 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_8_OAI21X1_112 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_51_5_1 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_16_DFFSR_271 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_6_NAND3X1_190 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_20_CLKBUF1_26 INVX1_1/gnd DFFSR_53/S FILL
XFILL_12_XOR2X1_6 BUFX2_99/A DFFSR_7/S FILL
XFILL_19_DFFSR_9 BUFX2_79/A DFFSR_6/S FILL
XFILL_19_CLKBUF1_29 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_43_DFFSR_93 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_8_DFFSR_158 INVX1_3/gnd DFFSR_23/S FILL
XFILL_49_DFFSR_189 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_18_CLKBUF1_32 DFFSR_1/gnd DFFSR_81/S FILL
XNAND3X1_226 INVX1_177/A NAND2X1_108/Y OAI21X1_79/Y OR2X2_3/gnd NAND3X1_226/Y DFFSR_60/S
+ NAND3X1
XFILL_4_AND2X2_2 BUFX2_99/A DFFSR_7/S FILL
XFILL_17_CLKBUF1_35 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_39_DFFSR_192 INVX1_1/gnd DFFSR_97/S FILL
XFILL_1_INVX1_135 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_27_DFFSR_43 BUFX2_98/A DFFSR_6/S FILL
XFILL_16_DFFSR_83 INVX1_3/gnd DFFSR_79/S FILL
XFILL_7_NAND3X1_124 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_2_DFFSR_268 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_16_CLKBUF1_38 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_29_DFFSR_195 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_11_DFFPOSX1_28 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_19_DFFSR_198 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_15_CLKBUF1_41 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_0_NAND2X1_105 OR2X2_6/gnd DFFSR_53/S FILL
XNOR2X1_80 NOR2X1_80/A NOR2X1_80/B NOR3X1_6/gnd NOR2X1_80/Y DFFSR_91/S NOR2X1
XFILL_14_CLKBUF1_44 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_13_CLKBUF1_47 BUFX2_98/A DFFSR_32/S FILL
XFILL_17_6_0 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_4_NOR2X1_77 INVX1_39/gnd DFFSR_34/S FILL
XFILL_40_DFFSR_5 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_21_DFFPOSX1_17 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_42_DFFSR_119 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_46_DFFSR_10 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_35_DFFSR_50 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_7_DFFSR_97 INVX1_1/gnd DFFSR_97/S FILL
XFILL_24_DFFSR_90 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_11_XNOR2X1_1 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_5_DFFSR_195 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_32_DFFSR_122 BUFX2_79/A DFFSR_7/S FILL
XFILL_46_DFFSR_226 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_5_NAND3X1_220 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_22_DFFSR_125 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_1_DFFPOSX1_39 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_36_DFFSR_229 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_1_AND2X2_39 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_12_DFFSR_128 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_6_BUFX2_35 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_26_DFFSR_232 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_2_AOI21X1_7 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_16_DFFSR_235 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_6_NAND3X1_154 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_43_DFFSR_57 BUFX2_79/A DFFSR_6/S FILL
XFILL_8_DFFSR_122 BUFX2_79/A DFFSR_7/S FILL
XFILL_32_DFFSR_97 INVX1_1/gnd DFFSR_97/S FILL
XFILL_4_INVX1_91 AND2X2_38/B DFFSR_23/S FILL
XFILL_49_DFFSR_153 INVX1_67/gnd DFFSR_201/S FILL
XNAND3X1_190 AOI21X1_26/C AOI21X1_26/B AOI21X1_26/A BUFX2_7/gnd NAND3X1_190/Y DFFSR_151/S
+ NAND3X1
XFILL_39_DFFSR_156 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_16_DFFSR_47 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_3_BUFX2_82 INVX1_1/gnd DFFSR_97/S FILL
XFILL_2_DFFSR_232 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_29_DFFSR_159 DFFSR_62/gnd DFFSR_208/S FILL
XNAND3X1_9 DFFSR_42/Q BUFX2_17/Y BUFX2_12/Y OR2X2_4/gnd NAND3X1_9/Y DFFSR_3/S NAND3X1
XFILL_43_DFFSR_263 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_19_DFFSR_162 BUFX2_99/A DFFSR_92/S FILL
XFILL_20_DFFPOSX1_47 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_33_DFFSR_266 INVX1_67/gnd DFFSR_201/S FILL
XFILL_27_1_0 INVX1_3/gnd DFFSR_79/S FILL
XNOR2X1_44 NOR2X1_44/A NOR2X1_44/B DFFSR_34/gnd NOR2X1_44/Y DFFSR_1/S NOR2X1
XFILL_4_NAND3X1_6 BUFX2_99/A DFFSR_92/S FILL
XFILL_23_DFFSR_269 INVX1_67/gnd DFFSR_201/S FILL
XFILL_13_CLKBUF1_11 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_4_NOR2X1_41 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_13_DFFSR_272 INVX1_3/gnd DFFSR_23/S FILL
XFILL_25_3_1 AND2X2_38/B DFFSR_23/S FILL
XFILL_12_CLKBUF1_14 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_7_OAI21X1_106 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_7_DFFSR_61 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_35_DFFSR_14 INVX1_1/gnd DFFSR_53/S FILL
XFILL_11_CLKBUF1_17 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_7_2_0 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_13_DFFSR_94 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_24_DFFSR_54 INVX1_39/gnd DFFSR_54/S FILL
XFILL_5_DFFSR_159 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_23_5_2 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_5_NAND3X1_184 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_10_CLKBUF1_20 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_46_DFFSR_190 INVX1_39/gnd DFFSR_34/S FILL
XFILL_9_DFFSR_266 INVX1_67/gnd DFFSR_201/S FILL
XFILL_36_DFFSR_193 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_5_4_1 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_26_DFFSR_196 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_9_CLKBUF1_23 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_7_DFFSR_8 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_8_CLKBUF1_26 INVX1_1/gnd DFFSR_53/S FILL
XFILL_16_DFFSR_199 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_3_6_2 INVX1_67/gnd DFFSR_175/S FILL
XFILL_6_NAND3X1_118 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_7_CLKBUF1_29 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_10_DFFPOSX1_22 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_32_DFFSR_61 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_4_INVX1_55 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_43_DFFSR_21 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_1_NOR2X1_78 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_6_CLKBUF1_32 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_49_DFFSR_117 BUFX2_77/gnd DFFSR_98/S FILL
XNAND3X1_154 INVX1_148/A NOR3X1_5/A INVX1_147/Y BUFX2_7/gnd INVX1_155/A DFFSR_216/S
+ NAND3X1
XFILL_5_CLKBUF1_35 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_39_DFFSR_120 INVX1_3/gnd DFFSR_23/S FILL
XCLKBUF1_32 BUFX2_3/Y DFFSR_1/gnd AOI21X1_3/B DFFSR_81/S CLKBUF1
XFILL_16_DFFSR_11 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_4_CLKBUF1_38 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_2_DFFSR_196 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_3_BUFX2_46 BUFX2_98/A DFFSR_6/S FILL
XFILL_29_DFFSR_123 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_43_DFFSR_227 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_3_CLKBUF1_41 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_8_AND2X2_37 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_20_DFFPOSX1_11 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_19_DFFSR_126 BUFX2_99/A DFFSR_7/S FILL
XFILL_33_DFFSR_230 INVX1_67/gnd DFFSR_201/S FILL
XFILL_2_CLKBUF1_44 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_23_DFFSR_233 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_1_CLKBUF1_47 BUFX2_98/A DFFSR_32/S FILL
XFILL_4_NAND3X1_214 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_40_DFFSR_68 BUFX2_98/A DFFSR_6/S FILL
XFILL_0_DFFPOSX1_33 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_13_DFFSR_236 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_33_0_2 INVX1_1/gnd DFFSR_53/S FILL
XFILL_7_DFFSR_25 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_13_DFFSR_58 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_5_DFFSR_123 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_24_DFFSR_18 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_0_BUFX2_93 AND2X2_38/B DFFSR_59/S FILL
XFILL_46_DFFSR_154 BUFX2_99/A DFFSR_7/S FILL
XFILL_5_NAND3X1_148 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_9_DFFSR_230 INVX1_67/gnd DFFSR_201/S FILL
XFILL_36_DFFSR_157 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_50_DFFSR_261 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_6_NOR2X1_6 BUFX2_98/A DFFSR_6/S FILL
XFILL_26_DFFSR_160 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_40_DFFSR_264 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_2_INVX1_207 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_48_DFFSR_75 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_16_DFFSR_163 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_30_DFFSR_267 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_1_NAND3X1_7 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_20_DFFSR_270 INVX1_39/gnd DFFSR_54/S FILL
XFILL_19_DFFPOSX1_41 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_4_DFFSR_72 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_32_DFFSR_25 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_21_DFFSR_65 BUFX2_79/A DFFSR_7/S FILL
XFILL_4_INVX1_19 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_1_NOR2X1_42 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_10_DFFSR_273 DFFSR_62/gnd DFFSR_208/S FILL
XNAND3X1_118 DFFSR_199/Q BUFX2_28/Y NOR2X1_31/Y DFFSR_62/gnd NAND3X1_118/Y DFFSR_62/S
+ NAND3X1
XFILL_3_NAND3X1_244 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_2_DFFSR_160 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_3_BUFX2_10 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_8_XOR2X1_2 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_43_DFFSR_191 INVX1_67/gnd DFFSR_175/S FILL
XFILL_6_OAI21X1_100 INVX1_3/gnd DFFSR_79/S FILL
XFILL_6_DFFSR_267 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_33_DFFSR_194 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_23_DFFSR_197 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_4_NAND3X1_178 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_1_CLKBUF1_11 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_1_INVX1_66 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_40_DFFSR_32 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_29_DFFSR_72 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_0_CLKBUF1_14 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_13_DFFSR_200 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_13_DFFSR_22 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_0_BUFX2_57 AND2X2_38/B DFFSR_23/S FILL
XFILL_46_DFFSR_118 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_5_NAND3X1_112 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_9_DFFSR_194 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_36_DFFSR_121 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_4_NOR3X1_3 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_50_DFFSR_225 INVX1_67/gnd DFFSR_175/S FILL
XFILL_18_DFFSR_6 BUFX2_79/A DFFSR_6/S FILL
XFILL_26_DFFSR_124 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_2_INVX1_171 BUFX2_98/A DFFSR_6/S FILL
XFILL_40_DFFSR_228 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_37_DFFSR_79 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_48_DFFSR_39 INVX1_3/gnd DFFSR_79/S FILL
XFILL_5_AND2X2_38 AND2X2_38/B DFFSR_59/S FILL
XFILL_16_DFFSR_127 BUFX2_99/A DFFSR_92/S FILL
XFILL_24_6_0 AND2X2_38/B DFFSR_59/S FILL
XFILL_30_DFFSR_231 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_6_AOI21X1_6 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_20_DFFSR_234 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_21_DFFSR_29 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_4_DFFSR_36 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_2_BUFX2_7 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_10_DFFSR_69 BUFX2_98/A DFFSR_32/S FILL
XFILL_10_DFFSR_237 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_3_NAND3X1_208 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_2_DFFSR_124 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_39_DFFSR_2 BUFX2_79/A DFFSR_7/S FILL
XFILL_43_DFFSR_155 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_45_DFFSR_86 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_6_DFFSR_231 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_33_DFFSR_158 INVX1_3/gnd DFFSR_23/S FILL
XFILL_47_DFFSR_262 BUFX2_98/A DFFSR_32/S FILL
XFILL_23_DFFSR_161 INVX1_67/gnd DFFSR_175/S FILL
XFILL_4_NAND3X1_142 INVX1_67/gnd DFFSR_175/S FILL
XFILL_37_DFFSR_265 INVX1_67/gnd DFFSR_175/S FILL
XFILL_1_INVX1_30 INVX1_1/gnd DFFSR_53/S FILL
XFILL_1_DFFSR_83 INVX1_3/gnd DFFSR_79/S FILL
XFILL_29_DFFSR_36 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_18_DFFSR_76 BUFX2_79/A DFFSR_7/S FILL
XFILL_24_DFFPOSX1_2 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_8_NAND3X1_5 BUFX2_99/A DFFSR_7/S FILL
XFILL_13_DFFSR_164 OR2X2_2/gnd DFFSR_216/S FILL
XOAI21X1_100 BUFX2_55/Y INVX1_197/Y NAND2X1_131/Y INVX1_3/gnd DFFSR_272/D DFFSR_79/S
+ OAI21X1
XFILL_9_DFFPOSX1_16 INVX1_67/gnd DFFSR_175/S FILL
XFILL_27_DFFSR_268 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_23_DFFPOSX1_5 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_6_NAND2X1_178 INVX1_1/gnd DFFSR_53/S FILL
XFILL_17_DFFSR_271 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_22_DFFPOSX1_8 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_0_BUFX2_21 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_9_DFFSR_158 INVX1_3/gnd DFFSR_23/S FILL
XFILL_18_DFFPOSX1_35 INVX1_39/gnd DFFSR_54/S FILL
XFILL_50_DFFSR_189 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_34_1_0 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_40_DFFSR_192 INVX1_1/gnd DFFSR_97/S FILL
XFILL_2_INVX1_135 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_9_DFFSR_90 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_37_DFFSR_43 BUFX2_98/A DFFSR_6/S FILL
XFILL_26_DFFSR_83 INVX1_3/gnd DFFSR_79/S FILL
XFILL_2_NAND3X1_238 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_3_DFFSR_268 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_30_DFFSR_195 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_32_3_1 INVX1_1/gnd DFFSR_97/S FILL
XFILL_20_DFFSR_198 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_10_DFFSR_33 BUFX2_98/A DFFSR_32/S FILL
XFILL_10_DFFSR_201 INVX1_67/gnd DFFSR_201/S FILL
XFILL_30_5_2 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_3_NAND3X1_172 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_5_NOR2X1_77 INVX1_39/gnd DFFSR_34/S FILL
XFILL_43_DFFSR_119 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_8_DFFPOSX1_46 INVX1_39/gnd DFFSR_34/S FILL
XFILL_45_DFFSR_50 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_34_DFFSR_90 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_12_XNOR2X1_1 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_6_DFFSR_195 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_33_DFFSR_122 BUFX2_79/A DFFSR_7/S FILL
XFILL_47_DFFSR_226 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_23_DFFSR_125 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_4_NAND3X1_106 INVX1_3/gnd DFFSR_23/S FILL
XFILL_1_DFFSR_47 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_37_DFFSR_229 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_18_DFFSR_40 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_2_AND2X2_39 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_5_BUFX2_75 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_13_DFFSR_128 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_27_DFFSR_232 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_6_NAND2X1_142 INVX1_67/gnd DFFSR_175/S FILL
XFILL_3_AOI21X1_7 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_17_DFFSR_235 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_6_DFFSR_5 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_9_DFFSR_122 BUFX2_79/A DFFSR_7/S FILL
XFILL_42_DFFSR_97 INVX1_1/gnd DFFSR_97/S FILL
XNAND2X1_178 XOR2X1_14/A XOR2X1_14/B INVX1_1/gnd NAND2X1_180/A DFFSR_53/S NAND2X1
XFILL_50_DFFSR_153 INVX1_67/gnd DFFSR_201/S FILL
XFILL_8_AOI21X1_70 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_3_AND2X2_6 BUFX2_99/A DFFSR_7/S FILL
XFILL_40_DFFSR_156 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_26_DFFSR_47 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_9_DFFSR_54 INVX1_39/gnd DFFSR_54/S FILL
XFILL_15_DFFSR_87 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_2_NAND3X1_202 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_3_DFFSR_232 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_30_DFFSR_159 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_44_DFFSR_263 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_20_DFFSR_162 BUFX2_99/A DFFSR_92/S FILL
XFILL_4_OR2X2_5 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_34_DFFSR_266 INVX1_67/gnd DFFSR_201/S FILL
XFILL_40_0_2 BUFX2_98/A DFFSR_6/S FILL
XFILL_5_NAND3X1_6 BUFX2_99/A DFFSR_92/S FILL
XFILL_10_DFFSR_165 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_24_DFFSR_269 INVX1_67/gnd DFFSR_201/S FILL
XFILL_3_NAND3X1_136 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_5_NOR2X1_41 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_30_DFFSR_9 BUFX2_79/A DFFSR_6/S FILL
XFILL_14_DFFSR_272 INVX1_3/gnd DFFSR_23/S FILL
XFILL_8_DFFPOSX1_10 INVX1_67/gnd DFFSR_201/S FILL
XFILL_45_DFFSR_14 INVX1_1/gnd DFFSR_53/S FILL
XFILL_5_NAND2X1_172 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_23_DFFSR_94 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_34_DFFSR_54 INVX1_39/gnd DFFSR_54/S FILL
XFILL_6_DFFSR_159 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_12_DFFPOSX1_2 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_47_DFFSR_190 INVX1_39/gnd DFFSR_34/S FILL
XFILL_11_DFFPOSX1_5 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_37_DFFSR_193 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_1_DFFSR_11 DFFSR_1/gnd DFFSR_1/S FILL
XBUFX2_79 BUFX2_79/A BUFX2_79/A BUFX2_79/Y DFFSR_7/S BUFX2
XFILL_0_DFFSR_269 INVX1_67/gnd DFFSR_201/S FILL
XFILL_5_BUFX2_39 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_10_DFFPOSX1_8 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_17_DFFPOSX1_29 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_27_DFFSR_196 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_6_NAND2X1_106 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_17_DFFSR_199 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_1_NAND3X1_232 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_3_INVX1_95 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_42_DFFSR_61 DFFSR_28/gnd DFFSR_8/S FILL
XNAND2X1_142 DFFPOSX1_37/Q INVX1_208/Y INVX1_67/gnd AOI21X1_47/A DFFSR_175/S NAND2X1
XFILL_2_NOR2X1_78 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_50_DFFSR_117 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_8_AOI21X1_34 INVX1_39/gnd DFFSR_34/S FILL
XFILL_27_DFFPOSX1_18 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_40_DFFSR_120 INVX1_3/gnd DFFSR_23/S FILL
XFILL_7_AOI21X1_37 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_9_DFFSR_18 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_26_DFFSR_11 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_15_DFFSR_51 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_2_NAND3X1_166 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_3_DFFSR_196 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_2_BUFX2_86 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_30_DFFSR_123 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_6_AOI21X1_40 INVX1_39/gnd DFFSR_54/S FILL
XFILL_44_DFFSR_227 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_20_DFFSR_126 BUFX2_99/A DFFSR_7/S FILL
XFILL_7_DFFPOSX1_40 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_34_DFFSR_230 INVX1_67/gnd DFFSR_201/S FILL
XFILL_5_AOI21X1_43 INVX1_3/gnd DFFSR_79/S FILL
XAOI21X1_40 AOI21X1_40/A AOI21X1_40/B INVX1_169/Y INVX1_39/gnd AOI21X1_40/Y DFFSR_54/S
+ AOI21X1
XFILL_10_DFFSR_129 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_4_AOI21X1_46 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_24_DFFSR_233 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_0_AOI21X1_8 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_50_DFFSR_68 BUFX2_98/A DFFSR_6/S FILL
XFILL_3_NAND3X1_100 AND2X2_38/B DFFSR_59/S FILL
XFILL_3_AOI21X1_49 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_20_2 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_14_DFFSR_236 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_2_AOI21X1_52 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_5_NAND2X1_136 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_6_DFFSR_65 BUFX2_79/A DFFSR_7/S FILL
XFILL_23_DFFSR_58 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_12_DFFSR_98 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_6_DFFSR_123 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_34_DFFSR_18 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_1_AOI21X1_55 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_47_DFFSR_154 BUFX2_99/A DFFSR_7/S FILL
XFILL_0_AOI21X1_58 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_31_6_0 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_37_DFFSR_157 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_51_DFFSR_261 BUFX2_77/gnd DFFSR_98/S FILL
XBUFX2_43 INVX1_59/Y AND2X2_38/B DFFSR_1/R DFFSR_23/S BUFX2
XFILL_0_DFFSR_233 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_27_DFFSR_160 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_3_OAI21X1_118 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_41_DFFSR_264 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_26_DFFPOSX1_48 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_3_INVX1_207 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_17_DFFSR_163 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_8_OAI21X1_82 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_17_DFFSR_3 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_1_NAND3X1_196 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_31_DFFSR_267 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_2_NAND3X1_7 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_7_OAI21X1_85 INVX1_39/gnd DFFSR_54/S FILL
XFILL_21_DFFSR_270 INVX1_39/gnd DFFSR_54/S FILL
XFILL_42_DFFSR_25 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_31_DFFSR_65 BUFX2_79/A DFFSR_7/S FILL
XFILL_3_INVX1_59 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_2_NOR2X1_42 BUFX2_8/gnd DFFSR_81/S FILL
XNAND2X1_106 BUFX2_56/Y DFFPOSX1_50/Q OR2X2_6/gnd XNOR2X1_2/B DFFSR_53/S NAND2X1
XFILL_6_OAI21X1_88 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_11_DFFSR_273 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_5_OAI21X1_91 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_1_BUFX2_4 OR2X2_6/gnd DFFSR_92/S FILL
XOAI21X1_88 DFFSR_260/S INVX1_184/Y OAI21X1_88/C DFFSR_5/gnd DFFSR_260/D DFFSR_5/S
+ OAI21X1
XFILL_15_DFFSR_15 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_2_NAND3X1_130 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_4_OAI21X1_94 INVX1_67/gnd DFFSR_175/S FILL
XFILL_3_DFFSR_160 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_2_BUFX2_50 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_44_DFFSR_191 INVX1_67/gnd DFFSR_175/S FILL
XFILL_3_OAI21X1_97 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_7_DFFSR_267 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_4_NAND2X1_166 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_34_DFFSR_194 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_4_AOI21X1_10 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_24_DFFSR_197 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_50_DFFSR_32 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_39_DFFSR_72 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_3_AOI21X1_13 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_14_DFFSR_200 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_2_AOI21X1_16 INVX1_67/gnd DFFSR_175/S FILL
XFILL_16_DFFPOSX1_23 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_6_DFFSR_29 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_41_1_0 BUFX2_98/A DFFSR_32/S FILL
XFILL_5_NAND2X1_100 INVX1_39/gnd DFFSR_54/S FILL
XFILL_23_DFFSR_22 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_0_DFFPOSX1_2 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_12_DFFSR_62 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_1_AOI21X1_19 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_47_DFFSR_118 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_0_NAND3X1_226 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_0_AOI21X1_22 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_39_3_1 BUFX2_79/A DFFSR_6/S FILL
XFILL_37_DFFSR_121 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_0_DFFSR_197 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_27_DFFSR_124 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_26_DFFPOSX1_12 AND2X2_38/B DFFSR_23/S FILL
XFILL_41_DFFSR_228 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_3_INVX1_171 BUFX2_98/A DFFSR_6/S FILL
XFILL_47_DFFSR_79 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_6_AND2X2_38 AND2X2_38/B DFFSR_59/S FILL
XFILL_17_DFFSR_127 BUFX2_99/A DFFSR_92/S FILL
XFILL_37_5_2 BUFX2_99/A DFFSR_7/S FILL
XFILL_8_OAI21X1_46 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_31_DFFSR_231 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_1_NAND3X1_160 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_7_AOI21X1_6 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_6_NAND2X1_67 AND2X2_38/B DFFSR_59/S FILL
XFILL_7_OAI21X1_49 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_21_DFFSR_234 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_31_DFFSR_29 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_3_DFFSR_76 BUFX2_79/A DFFSR_7/S FILL
XFILL_3_INVX1_23 BUFX2_99/A DFFSR_7/S FILL
XFILL_6_DFFPOSX1_34 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_20_DFFSR_69 BUFX2_98/A DFFSR_32/S FILL
XFILL_5_NAND2X1_70 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_6_OAI21X1_52 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_11_DFFSR_237 DFFSR_1/gnd DFFSR_1/S FILL
XNAND2X1_67 AND2X2_35/A INVX1_175/A AND2X2_38/B INVX1_144/A DFFSR_59/S NAND2X1
XFILL_4_NAND2X1_73 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_5_OAI21X1_55 DFFSR_62/gnd DFFSR_208/S FILL
XOAI21X1_52 OAI21X1_54/A OAI21X1_54/B OAI21X1_53/C XOR2X1_1/gnd OAI21X1_52/Y DFFSR_208/S
+ OAI21X1
XFILL_42_2 BUFX2_98/A DFFSR_32/S FILL
XFILL_3_NAND2X1_76 INVX1_3/gnd DFFSR_23/S FILL
XFILL_3_DFFSR_124 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_4_OAI21X1_58 INVX1_39/gnd DFFSR_54/S FILL
XFILL_2_BUFX2_14 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_7_XOR2X1_6 BUFX2_99/A DFFSR_7/S FILL
XFILL_44_DFFSR_155 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_10_AOI22X1_2 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_3_OAI21X1_61 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_2_NAND2X1_79 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_7_DFFSR_231 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_34_DFFSR_158 INVX1_3/gnd DFFSR_23/S FILL
XFILL_4_NAND2X1_130 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_1_NAND2X1_82 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_48_DFFSR_262 BUFX2_98/A DFFSR_32/S FILL
XFILL_2_OAI21X1_64 INVX1_1/gnd DFFSR_53/S FILL
XFILL_24_DFFSR_161 INVX1_67/gnd DFFSR_175/S FILL
XFILL_38_DFFSR_265 INVX1_67/gnd DFFSR_175/S FILL
XFILL_1_OAI21X1_67 INVX1_1/gnd DFFSR_97/S FILL
XFILL_0_NAND2X1_85 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_39_DFFSR_36 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_28_DFFSR_76 BUFX2_79/A DFFSR_7/S FILL
XFILL_0_INVX1_70 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_0_INVX1_208 INVX1_39/gnd DFFSR_34/S FILL
XFILL_14_DFFSR_164 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_0_OAI21X1_70 INVX1_3/gnd DFFSR_23/S FILL
XFILL_28_DFFSR_268 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_2_OAI21X1_112 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_18_DFFSR_271 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_25_DFFPOSX1_42 INVX1_39/gnd DFFSR_34/S FILL
XFILL_12_DFFSR_26 BUFX2_79/A DFFSR_6/S FILL
XFILL_0_NAND3X1_190 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_9_NAND3X1_245 OR2X2_4/gnd DFFSR_3/S FILL
XDFFSR_6 DFFSR_6/Q DFFSR_2/CLK DFFSR_2/R DFFSR_6/S DFFSR_6/D BUFX2_79/A DFFSR_6/S
+ DFFSR
XFILL_5_DFFSR_2 BUFX2_79/A DFFSR_7/S FILL
XFILL_0_DFFSR_161 INVX1_67/gnd DFFSR_175/S FILL
XFILL_47_0_2 DFFSR_8/gnd DFFSR_60/S FILL
XDFFSR_271 INVX1_196/A CLKBUF1_48/Y DFFSR_266/R DFFSR_81/S DFFSR_271/D BUFX2_8/gnd
+ DFFSR_81/S DFFSR
XFILL_41_DFFSR_192 INVX1_1/gnd DFFSR_97/S FILL
XFILL_47_DFFSR_43 BUFX2_98/A DFFSR_6/S FILL
XFILL_3_INVX1_135 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_36_DFFSR_83 INVX1_3/gnd DFFSR_79/S FILL
XFILL_4_DFFSR_268 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_8_OAI21X1_10 BUFX2_79/A DFFSR_7/S FILL
XFILL_31_DFFSR_195 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_1_NAND3X1_124 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_6_NAND2X1_31 INVX1_3/gnd DFFSR_23/S FILL
XFILL_7_OAI21X1_13 INVX1_39/gnd DFFSR_54/S FILL
XFILL_21_DFFSR_198 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_3_DFFSR_40 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_20_DFFSR_33 BUFX2_98/A DFFSR_32/S FILL
XFILL_6_OAI21X1_16 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_5_NAND2X1_34 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_11_DFFSR_201 INVX1_67/gnd DFFSR_201/S FILL
XFILL_3_NAND2X1_160 NOR3X1_6/gnd DFFSR_79/S FILL
XNAND2X1_31 AND2X2_18/B AND2X2_15/Y INVX1_3/gnd OAI22X1_45/D DFFSR_23/S NAND2X1
XFILL_3_OR2X2_2 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_4_NAND2X1_37 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_5_OAI21X1_19 BUFX2_98/A DFFSR_32/S FILL
XFILL_6_NOR2X1_77 INVX1_39/gnd DFFSR_34/S FILL
XOAI21X1_16 INVX1_117/Y OAI21X1_9/B OAI21X1_16/C XOR2X1_4/gnd NOR2X1_57/B DFFSR_97/S
+ OAI21X1
XFILL_3_NAND2X1_40 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_4_OAI21X1_22 DFFSR_34/gnd DFFSR_34/S FILL
XDFFPOSX1_34 DFFPOSX1_34/Q CLKBUF1_43/Y AOI21X1_49/Y OR2X2_2/gnd DFFSR_216/S DFFPOSX1
XFILL_13_XOR2X1_3 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_44_DFFSR_119 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_29_DFFSR_6 BUFX2_79/A DFFSR_6/S FILL
XFILL_15_DFFPOSX1_17 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_2_NAND2X1_43 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_3_OAI21X1_25 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_44_DFFSR_90 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_13_XNOR2X1_1 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_7_DFFSR_195 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_34_DFFSR_122 BUFX2_79/A DFFSR_7/S FILL
XFILL_1_NAND2X1_46 INVX1_39/gnd DFFSR_34/S FILL
XFILL_2_OAI21X1_28 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_48_DFFSR_226 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_24_DFFSR_125 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_13_1_1 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_0_NAND2X1_49 INVX1_3/gnd DFFSR_79/S FILL
XFILL_1_OAI21X1_31 AND2X2_38/B DFFSR_23/S FILL
XFILL_38_DFFSR_229 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_28_DFFSR_40 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_0_INVX1_172 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_17_DFFSR_80 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_0_DFFSR_87 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_0_INVX1_34 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_3_AND2X2_39 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_14_DFFSR_128 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_0_OAI21X1_34 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_28_DFFSR_232 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_4_AOI21X1_7 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_11_3_2 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_18_DFFSR_235 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_0_NAND3X1_154 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_50_DFFSR_2 BUFX2_79/A DFFSR_7/S FILL
XFILL_5_DFFPOSX1_28 BUFX2_72/gnd DFFSR_201/S FILL
XDFFSR_235 DFFSR_235/Q CLKBUF1_2/Y BUFX2_67/Y DFFSR_216/S DFFSR_235/D OR2X2_2/gnd
+ DFFSR_216/S DFFSR
XFILL_0_DFFSR_125 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_41_DFFSR_156 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_36_DFFSR_47 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_8_DFFSR_94 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_25_DFFSR_87 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_4_DFFSR_232 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_5_AOI22X1_12 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_31_DFFSR_159 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_45_DFFSR_263 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_4_AOI22X1_15 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_21_DFFSR_162 BUFX2_99/A DFFSR_92/S FILL
XFILL_14_DFFPOSX1_47 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_35_DFFSR_266 INVX1_67/gnd DFFSR_201/S FILL
XFILL_3_AOI22X1_18 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_6_NAND3X1_6 BUFX2_99/A DFFSR_92/S FILL
XFILL_11_DFFSR_165 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_3_NAND2X1_124 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_25_DFFSR_269 INVX1_67/gnd DFFSR_201/S FILL
XINVX1_8 INVX1_8/A OR2X2_4/gnd INVX1_8/Y DFFSR_3/S INVX1
XFILL_2_AOI22X1_21 AND2X2_38/B DFFSR_59/S FILL
XFILL_6_NOR2X1_41 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_38_6_0 BUFX2_79/A DFFSR_7/S FILL
XFILL_15_DFFSR_272 INVX1_3/gnd DFFSR_23/S FILL
XFILL_11_OAI22X1_42 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_1_AOI22X1_24 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_10_OAI22X1_45 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_0_AOI22X1_27 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_33_DFFSR_94 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_44_DFFSR_54 INVX1_39/gnd DFFSR_54/S FILL
XFILL_1_OAI21X1_106 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_7_DFFSR_159 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_24_DFFPOSX1_36 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_9_NAND3X1_63 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_1_NAND2X1_10 BUFX2_79/A DFFSR_7/S FILL
XFILL_48_DFFSR_190 INVX1_39/gnd DFFSR_34/S FILL
XAND2X2_3 INVX1_3/A NOR3X1_1/A INVX1_1/gnd AND2X2_3/Y DFFSR_53/S AND2X2
XFILL_8_NAND3X1_66 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_9_OAI22X1_48 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_38_DFFSR_193 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_0_NAND2X1_13 BUFX2_99/A DFFSR_92/S FILL
XFILL_0_INVX1_136 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_8_NAND3X1_239 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_17_DFFSR_44 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_0_DFFSR_51 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_1_DFFSR_269 INVX1_67/gnd DFFSR_201/S FILL
XFILL_7_NAND3X1_69 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_8_OAI22X1_51 INVX1_39/gnd DFFSR_54/S FILL
XFILL_4_BUFX2_79 BUFX2_79/A DFFSR_7/S FILL
XFILL_28_DFFSR_196 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_6_NAND3X1_72 INVX1_39/gnd DFFSR_34/S FILL
XFILL_18_DFFSR_199 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_5_NAND3X1_75 BUFX2_79/A DFFSR_7/S FILL
XFILL_0_NAND3X1_118 DFFSR_62/gnd DFFSR_62/S FILL
XNAND3X1_72 NOR2X1_32/Y NOR2X1_35/Y NOR2X1_37/Y INVX1_39/gnd NAND3X1_72/Y DFFSR_34/S
+ NAND3X1
XFILL_9_NAND3X1_173 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_4_NAND3X1_78 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_3_NOR2X1_78 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_51_DFFSR_117 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_3_NAND3X1_81 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_2_NAND2X1_154 OR2X2_4/gnd DFFSR_3/S FILL
XDFFSR_199 DFFSR_199/Q CLKBUF1_20/Y BUFX2_66/Y DFFSR_208/S DFFSR_143/Q XOR2X1_1/gnd
+ DFFSR_208/S DFFSR
XFILL_41_DFFSR_120 INVX1_3/gnd DFFSR_23/S FILL
XFILL_2_NAND3X1_84 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_8_DFFSR_58 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_36_DFFSR_11 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_14_DFFSR_91 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_25_DFFSR_51 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_4_DFFSR_196 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_10_XNOR2X1_2 BUFX2_98/A DFFSR_6/S FILL
XFILL_31_DFFSR_123 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_1_NAND3X1_87 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_45_DFFSR_227 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_0_BUFX2_1 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_21_DFFSR_126 BUFX2_99/A DFFSR_7/S FILL
XFILL_0_NAND3X1_90 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_35_DFFSR_230 INVX1_67/gnd DFFSR_201/S FILL
XFILL_14_DFFPOSX1_11 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_48_1_0 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_0_AND2X2_40 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_11_DFFSR_129 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_25_DFFSR_233 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_1_AOI21X1_8 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_15_DFFSR_236 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_46_3_1 DFFSR_8/gnd DFFSR_8/S FILL
XINVX1_92 INVX1_92/A AND2X2_38/B INVX1_92/Y DFFSR_23/S INVX1
XFILL_33_DFFSR_58 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_22_DFFSR_98 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_44_DFFSR_18 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_7_DFFSR_123 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_9_NAND3X1_27 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_48_DFFSR_154 BUFX2_99/A DFFSR_7/S FILL
XFILL_44_5_2 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_9_OAI22X1_12 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_8_NAND3X1_30 BUFX2_79/A DFFSR_6/S FILL
XFILL_38_DFFSR_157 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_0_INVX1_100 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_0_DFFSR_15 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_8_NAND3X1_203 INVX1_1/gnd DFFSR_97/S FILL
XINVX1_210 INVX1_3/A NOR3X1_6/gnd NOR3X1_6/B DFFSR_79/S INVX1
XFILL_1_DFFSR_233 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_8_OAI22X1_15 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_7_NAND3X1_33 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_4_BUFX2_43 AND2X2_38/B DFFSR_23/S FILL
XFILL_28_DFFSR_160 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_4_DFFPOSX1_22 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_42_DFFSR_264 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_7_OAI22X1_18 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_6_NAND3X1_36 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_4_INVX1_207 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_18_DFFSR_163 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_32_DFFSR_267 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_5_NAND3X1_39 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_6_OAI22X1_21 BUFX2_98/A DFFSR_32/S FILL
XFILL_41_DFFSR_9 BUFX2_79/A DFFSR_6/S FILL
XFILL_3_NAND3X1_7 OR2X2_6/gnd DFFSR_92/S FILL
XNAND3X1_36 NAND3X1_36/A NAND3X1_33/Y AND2X2_10/Y DFFSR_8/gnd NOR2X1_20/A DFFSR_8/S
+ NAND3X1
XFILL_22_DFFSR_270 INVX1_39/gnd DFFSR_54/S FILL
XFILL_9_NAND3X1_137 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_5_OAI22X1_24 BUFX2_98/A DFFSR_32/S FILL
XFILL_4_NAND3X1_42 BUFX2_79/A DFFSR_6/S FILL
XFILL_41_DFFSR_65 BUFX2_79/A DFFSR_7/S FILL
XFILL_2_INVX1_99 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_3_NOR2X1_42 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_13_DFFPOSX1_41 DFFSR_8/gnd DFFSR_60/S FILL
XOAI22X1_21 INVX1_49/Y OAI22X1_6/B INVX1_50/Y OAI22X1_6/D BUFX2_98/A NOR2X1_25/A DFFSR_32/S
+ OAI22X1
XFILL_12_DFFSR_273 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_4_OAI22X1_27 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_3_NAND3X1_45 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_2_NAND2X1_118 NOR3X1_6/gnd DFFSR_79/S FILL
XDFFSR_163 DFFSR_163/Q CLKBUF1_29/Y BUFX2_66/Y DFFSR_1/S INVX1_80/A DFFSR_1/gnd DFFSR_1/S
+ DFFSR
XFILL_12_4_0 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_2_NAND3X1_48 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_3_OAI22X1_30 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_8_DFFSR_22 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_25_DFFSR_15 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_14_DFFSR_55 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_4_DFFSR_160 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_1_BUFX2_90 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_1_NAND3X1_51 BUFX2_99/A DFFSR_7/S FILL
XFILL_2_OAI22X1_33 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_45_DFFSR_191 INVX1_67/gnd DFFSR_175/S FILL
XFILL_10_6_1 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_1_OAI22X1_36 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_0_NAND3X1_54 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_8_DFFSR_267 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_35_DFFSR_194 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_0_OAI21X1_100 INVX1_3/gnd DFFSR_79/S FILL
XFILL_23_DFFPOSX1_30 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_0_OAI22X1_39 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_25_DFFSR_197 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_49_DFFSR_72 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_7_3 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_7_NAND3X1_233 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_15_DFFSR_200 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_54_0_2 DFFSR_5/gnd DFFSR_5/S FILL
XINVX1_56 DFFSR_24/Q BUFX2_98/A INVX1_56/Y DFFSR_6/S INVX1
XFILL_33_DFFSR_22 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_5_DFFSR_69 BUFX2_98/A DFFSR_32/S FILL
XFILL_22_DFFSR_62 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_0_NOR2X1_79 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_48_DFFSR_118 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_38_DFFSR_121 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_8_NAND3X1_167 XOR2X1_1/gnd DFFSR_208/S FILL
XINVX1_174 INVX1_174/A OR2X2_4/gnd OR2X2_3/B DFFSR_3/S INVX1
XFILL_1_DFFSR_197 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_28_DFFSR_124 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_1_NAND2X1_148 INVX1_67/gnd DFFSR_175/S FILL
XFILL_42_DFFSR_228 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_4_INVX1_171 BUFX2_98/A DFFSR_6/S FILL
XFILL_7_AND2X2_38 AND2X2_38/B DFFSR_59/S FILL
XFILL_18_DFFSR_127 BUFX2_99/A DFFSR_92/S FILL
XFILL_32_DFFSR_231 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_8_AOI21X1_6 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_22_DFFSR_234 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_2_INVX1_63 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_41_DFFSR_29 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_30_DFFSR_69 BUFX2_98/A DFFSR_32/S FILL
XFILL_12_DFFSR_237 DFFSR_1/gnd DFFSR_1/S FILL
XDFFSR_127 BUFX2_88/A CLKBUF1_5/Y DFFSR_7/R DFFSR_92/S INVX1_51/A BUFX2_99/A DFFSR_92/S
+ DFFSR
XFILL_2_NAND3X1_12 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_20_1_1 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_14_DFFSR_19 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_4_DFFSR_124 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_1_BUFX2_54 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_1_NAND3X1_15 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_2_0_0 INVX1_67/gnd DFFSR_201/S FILL
XFILL_45_DFFSR_155 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_11_AOI22X1_2 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_0_NAND3X1_18 BUFX2_79/A DFFSR_7/S FILL
XFILL_8_DFFSR_231 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_35_DFFSR_158 INVX1_3/gnd DFFSR_23/S FILL
XFILL_18_3_2 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_49_DFFSR_262 BUFX2_98/A DFFSR_32/S FILL
XFILL_28_DFFSR_3 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_0_2_1 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_25_DFFSR_161 INVX1_67/gnd DFFSR_175/S FILL
XFILL_39_DFFSR_265 INVX1_67/gnd DFFSR_175/S FILL
XFILL_49_DFFSR_36 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_38_DFFSR_76 BUFX2_79/A DFFSR_7/S FILL
XFILL_1_INVX1_208 INVX1_39/gnd DFFSR_34/S FILL
XFILL_15_DFFSR_164 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_7_NAND3X1_197 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_29_DFFSR_268 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_0_NAND3X1_8 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_3_DFFPOSX1_16 INVX1_67/gnd DFFSR_175/S FILL
XFILL_0_NAND2X1_178 INVX1_1/gnd DFFSR_53/S FILL
XINVX1_20 DFFSR_75/Q NOR3X1_6/gnd INVX1_20/Y DFFSR_79/S INVX1
XDFFSR_73 INVX1_6/A CLKBUF1_18/Y DFFSR_73/R DFFSR_51/S DFFSR_73/D OR2X2_1/gnd DFFSR_51/S
+ DFFSR
XFILL_19_DFFSR_271 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_5_DFFSR_33 BUFX2_98/A DFFSR_32/S FILL
XFILL_22_DFFSR_26 BUFX2_79/A DFFSR_6/S FILL
XFILL_11_DFFSR_66 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_0_NOR2X1_43 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_8_NAND3X1_131 AND2X2_38/B DFFSR_59/S FILL
XINVX1_138 INVX1_138/A DFFSR_1/gnd AOI21X1_8/A DFFSR_81/S INVX1
XFILL_1_DFFSR_161 INVX1_67/gnd DFFSR_175/S FILL
XFILL_12_DFFPOSX1_35 INVX1_39/gnd DFFSR_54/S FILL
XFILL_1_NAND2X1_112 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_42_DFFSR_192 INVX1_1/gnd DFFSR_97/S FILL
XFILL_46_DFFSR_83 INVX1_3/gnd DFFSR_79/S FILL
XFILL_5_DFFSR_268 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_32_DFFSR_195 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_45_6_0 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_22_DFFSR_198 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_2_INVX1_27 BUFX2_99/A DFFSR_7/S FILL
XFILL_2_DFFSR_80 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_30_DFFSR_33 BUFX2_98/A DFFSR_32/S FILL
XFILL_19_DFFSR_73 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_12_DFFSR_201 INVX1_67/gnd DFFSR_201/S FILL
XFILL_22_DFFPOSX1_24 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_6_NAND3X1_227 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_1_BUFX2_18 BUFX2_98/A DFFSR_32/S FILL
XFILL_4_INVX1_1 INVX1_1/gnd DFFSR_53/S FILL
XFILL_45_DFFSR_119 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_2_DFFPOSX1_46 INVX1_39/gnd DFFSR_34/S FILL
XFILL_14_XNOR2X1_1 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_8_DFFSR_195 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_35_DFFSR_122 BUFX2_79/A DFFSR_7/S FILL
XNOR3X1_4 NOR3X1_4/A NOR3X1_4/B NOR3X1_4/C NOR3X1_6/gnd NOR3X1_4/Y DFFSR_91/S NOR3X1
XFILL_49_DFFSR_226 DFFSR_4/gnd DFFSR_98/S FILL
XAND2X2_42 XOR2X1_10/A XOR2X1_10/B INVX1_3/gnd AND2X2_42/Y DFFSR_23/S AND2X2
XFILL_25_DFFSR_125 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_39_DFFSR_229 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_38_DFFSR_40 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_1_INVX1_172 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_27_DFFSR_80 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_4_AND2X2_39 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_15_DFFSR_128 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_7_NAND3X1_161 AND2X2_38/B DFFSR_23/S FILL
XFILL_29_DFFSR_232 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_5_AOI21X1_7 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_0_NAND2X1_142 INVX1_67/gnd DFFSR_175/S FILL
XFILL_19_DFFSR_235 OR2X2_2/gnd DFFSR_216/S FILL
XDFFSR_37 DFFSR_45/D DFFSR_85/CLK DFFSR_3/R DFFSR_60/S INVX1_35/A DFFSR_8/gnd DFFSR_60/S
+ DFFSR
XFILL_11_DFFSR_30 BUFX2_98/A DFFSR_32/S FILL
XINVX1_102 INVX1_102/A OR2X2_1/gnd INVX1_102/Y DFFSR_59/S INVX1
XFILL_1_DFFSR_125 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_42_DFFSR_156 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_51_4 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_35_DFFSR_87 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_46_DFFSR_47 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_5_DFFSR_232 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_32_DFFSR_159 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_46_DFFSR_263 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_53_3_1 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_22_DFFSR_162 BUFX2_99/A DFFSR_92/S FILL
XFILL_2_DFFSR_44 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_36_DFFSR_266 INVX1_67/gnd DFFSR_201/S FILL
XFILL_19_DFFSR_37 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_7_NAND3X1_6 BUFX2_99/A DFFSR_92/S FILL
XFILL_12_DFFSR_165 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_6_BUFX2_72 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_26_DFFSR_269 INVX1_67/gnd DFFSR_201/S FILL
XFILL_8_OAI21X1_113 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_51_5_2 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_16_DFFSR_272 INVX1_3/gnd DFFSR_23/S FILL
XFILL_6_NAND3X1_191 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_20_CLKBUF1_27 INVX1_1/gnd DFFSR_97/S FILL
XFILL_12_XOR2X1_7 BUFX2_98/A DFFSR_6/S FILL
XFILL_2_DFFPOSX1_10 INVX1_67/gnd DFFSR_201/S FILL
XFILL_19_CLKBUF1_30 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_43_DFFSR_94 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_8_DFFSR_159 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_18_CLKBUF1_33 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_49_DFFSR_190 INVX1_39/gnd DFFSR_34/S FILL
XNAND3X1_227 NAND3X1_227/A NAND3X1_226/Y INVX1_178/Y DFFSR_4/gnd NAND3X1_235/C DFFSR_4/S
+ NAND3X1
XFILL_39_DFFSR_193 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_4_AND2X2_3 INVX1_1/gnd DFFSR_53/S FILL
XFILL_17_CLKBUF1_36 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_1_INVX1_136 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_27_DFFSR_44 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_16_DFFSR_84 BUFX2_99/A DFFSR_7/S FILL
XFILL_2_DFFSR_269 INVX1_67/gnd DFFSR_201/S FILL
XFILL_7_NAND3X1_125 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_29_DFFSR_196 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_16_CLKBUF1_39 INVX1_1/gnd DFFSR_53/S FILL
XFILL_11_DFFPOSX1_29 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_15_CLKBUF1_42 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_0_NAND2X1_106 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_19_4_0 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_19_DFFSR_199 XOR2X1_1/gnd DFFSR_208/S FILL
XNOR2X1_81 NOR2X1_81/A NOR2X1_81/B XOR2X1_4/gnd NOR2X1_81/Y DFFSR_97/S NOR2X1
XFILL_14_CLKBUF1_45 BUFX2_79/A DFFSR_7/S FILL
XFILL_40_DFFSR_6 BUFX2_79/A DFFSR_6/S FILL
XFILL_4_NOR2X1_78 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_13_CLKBUF1_48 INVX1_3/gnd DFFSR_79/S FILL
XFILL_17_6_1 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_42_DFFSR_120 INVX1_3/gnd DFFSR_23/S FILL
XFILL_21_DFFPOSX1_18 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_7_DFFSR_98 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_24_DFFSR_91 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_35_DFFSR_51 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_46_DFFSR_11 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_5_DFFSR_196 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_11_XNOR2X1_2 BUFX2_98/A DFFSR_6/S FILL
XFILL_32_DFFSR_123 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_46_DFFSR_227 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_5_NAND3X1_221 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_22_DFFSR_126 BUFX2_99/A DFFSR_7/S FILL
XFILL_36_DFFSR_230 INVX1_67/gnd DFFSR_201/S FILL
XFILL_1_DFFPOSX1_40 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_1_AND2X2_40 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_6_BUFX2_36 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_12_DFFSR_129 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_26_DFFSR_233 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_11_1 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_2_AOI21X1_8 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_16_DFFSR_236 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_6_NAND3X1_155 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_43_DFFSR_58 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_4_INVX1_92 AND2X2_38/B DFFSR_23/S FILL
XFILL_32_DFFSR_98 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_8_DFFSR_123 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_49_DFFSR_154 BUFX2_99/A DFFSR_7/S FILL
XNAND3X1_191 NOR3X1_5/Y NAND3X1_187/Y NAND3X1_190/Y BUFX2_7/gnd NAND2X1_90/A DFFSR_151/S
+ NAND3X1
XFILL_39_DFFSR_157 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_1_INVX1_100 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_16_DFFSR_48 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_2_DFFSR_233 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_3_BUFX2_83 BUFX2_79/A DFFSR_7/S FILL
XFILL_29_DFFSR_160 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_43_DFFSR_264 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_20_DFFPOSX1_48 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_19_DFFSR_163 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_33_DFFSR_267 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_4_NAND3X1_7 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_27_1_1 INVX1_3/gnd DFFSR_79/S FILL
XNOR2X1_45 NOR2X1_45/A NOR2X1_45/B DFFSR_34/gnd NOR2X1_45/Y DFFSR_1/S NOR2X1
XFILL_23_DFFSR_270 INVX1_39/gnd DFFSR_54/S FILL
XFILL_9_0_0 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_13_CLKBUF1_12 AND2X2_38/B DFFSR_23/S FILL
XFILL_4_NOR2X1_42 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_13_DFFSR_273 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_25_3_2 AND2X2_38/B DFFSR_23/S FILL
XFILL_12_CLKBUF1_15 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_7_OAI21X1_107 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_7_2_1 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_35_DFFSR_15 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_24_DFFSR_55 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_11_CLKBUF1_18 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_7_DFFSR_62 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_13_DFFSR_95 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_5_DFFSR_160 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_46_DFFSR_191 INVX1_67/gnd DFFSR_175/S FILL
XFILL_10_CLKBUF1_21 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_5_NAND3X1_185 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_9_DFFSR_267 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_5_4_2 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_36_DFFSR_194 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_9_CLKBUF1_24 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_26_DFFSR_197 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_7_DFFSR_9 BUFX2_79/A DFFSR_6/S FILL
XFILL_16_DFFSR_200 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_8_CLKBUF1_27 INVX1_1/gnd DFFSR_97/S FILL
XFILL_6_NAND3X1_119 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_7_CLKBUF1_30 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_10_DFFPOSX1_23 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_43_DFFSR_22 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_4_INVX1_56 BUFX2_98/A DFFSR_6/S FILL
XFILL_32_DFFSR_62 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_6_CLKBUF1_33 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_1_NOR2X1_79 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_49_DFFSR_118 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_5_CLKBUF1_36 NOR3X1_6/gnd DFFSR_79/S FILL
XNAND3X1_155 BUFX2_54/Y NOR3X1_5/A INVX1_147/Y BUFX2_7/gnd OAI21X1_35/C DFFSR_216/S
+ NAND3X1
XFILL_52_6_0 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_39_DFFSR_121 OR2X2_6/gnd DFFSR_53/S FILL
XCLKBUF1_33 BUFX2_4/Y XOR2X1_4/gnd DFFSR_79/CLK DFFSR_91/S CLKBUF1
XFILL_16_DFFSR_12 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_4_CLKBUF1_39 INVX1_1/gnd DFFSR_53/S FILL
XFILL_2_DFFSR_197 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_3_BUFX2_47 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_29_DFFSR_124 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_3_CLKBUF1_42 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_43_DFFSR_228 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_20_DFFPOSX1_12 AND2X2_38/B DFFSR_23/S FILL
XFILL_8_AND2X2_38 AND2X2_38/B DFFSR_59/S FILL
XFILL_19_DFFSR_127 BUFX2_99/A DFFSR_92/S FILL
XFILL_2_CLKBUF1_45 BUFX2_79/A DFFSR_7/S FILL
XFILL_33_DFFSR_231 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_9_AOI21X1_6 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_23_DFFSR_234 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_1_CLKBUF1_48 INVX1_3/gnd DFFSR_79/S FILL
XFILL_4_NAND3X1_215 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_40_DFFSR_69 BUFX2_98/A DFFSR_32/S FILL
XFILL_13_DFFSR_237 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_0_DFFPOSX1_34 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_33_1 INVX1_1/gnd DFFSR_97/S FILL
XFILL_24_DFFSR_19 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_7_DFFSR_26 BUFX2_79/A DFFSR_6/S FILL
XFILL_13_DFFSR_59 AND2X2_38/B DFFSR_59/S FILL
XFILL_5_DFFSR_124 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_0_BUFX2_94 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_46_DFFSR_155 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_5_NAND3X1_149 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_9_DFFSR_231 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_36_DFFSR_158 INVX1_3/gnd DFFSR_23/S FILL
XFILL_50_DFFSR_262 BUFX2_98/A DFFSR_32/S FILL
XFILL_6_NOR2X1_7 BUFX2_98/A DFFSR_32/S FILL
XFILL_26_DFFSR_161 INVX1_67/gnd DFFSR_175/S FILL
XFILL_40_DFFSR_265 INVX1_67/gnd DFFSR_175/S FILL
XFILL_48_DFFSR_76 BUFX2_79/A DFFSR_7/S FILL
XFILL_2_INVX1_208 INVX1_39/gnd DFFSR_34/S FILL
XFILL_16_DFFSR_164 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_30_DFFSR_268 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_1_NAND3X1_8 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_20_DFFSR_271 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_4_DFFSR_73 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_21_DFFSR_66 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_32_DFFSR_26 BUFX2_79/A DFFSR_6/S FILL
XFILL_19_DFFPOSX1_42 INVX1_39/gnd DFFSR_34/S FILL
XFILL_1_NOR2X1_43 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_10_DFFSR_274 BUFX2_72/gnd DFFSR_276/S FILL
XNAND3X1_119 NAND3X1_117/Y NAND3X1_118/Y AOI22X1_15/Y DFFSR_46/gnd NOR2X1_55/B DFFSR_54/S
+ NAND3X1
XFILL_3_NAND3X1_245 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_2_DFFSR_161 INVX1_67/gnd DFFSR_175/S FILL
XFILL_3_BUFX2_11 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_8_XOR2X1_3 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_43_DFFSR_192 INVX1_1/gnd DFFSR_97/S FILL
XFILL_6_DFFSR_268 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_6_OAI21X1_101 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_33_DFFSR_195 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_23_DFFSR_198 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_4_NAND3X1_179 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_1_CLKBUF1_12 AND2X2_38/B DFFSR_23/S FILL
XFILL_1_INVX1_67 INVX1_67/gnd DFFSR_201/S FILL
XFILL_40_DFFSR_33 BUFX2_98/A DFFSR_32/S FILL
XFILL_29_DFFSR_73 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_13_DFFSR_201 INVX1_67/gnd DFFSR_201/S FILL
XFILL_0_CLKBUF1_15 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_13_DFFSR_23 AND2X2_38/B DFFSR_23/S FILL
XFILL_0_BUFX2_58 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_46_DFFSR_119 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_5_NAND3X1_113 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_15_XNOR2X1_1 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_9_DFFSR_195 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_36_DFFSR_122 BUFX2_79/A DFFSR_7/S FILL
XFILL_4_NOR3X1_4 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_50_DFFSR_226 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_26_4_0 INVX1_3/gnd DFFSR_23/S FILL
XFILL_18_DFFSR_7 BUFX2_79/A DFFSR_7/S FILL
XFILL_26_DFFSR_125 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_48_DFFSR_40 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_2_INVX1_172 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_40_DFFSR_229 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_37_DFFSR_80 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_5_AND2X2_39 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_16_DFFSR_128 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_24_6_1 AND2X2_38/B DFFSR_59/S FILL
XFILL_30_DFFSR_232 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_6_AOI21X1_7 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_20_DFFSR_235 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_6_5_0 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_4_DFFSR_37 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_10_DFFSR_70 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_21_DFFSR_30 BUFX2_98/A DFFSR_32/S FILL
XFILL_2_BUFX2_8 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_10_DFFSR_238 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_3_NAND3X1_209 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_2_DFFSR_125 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_43_DFFSR_156 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_55_1 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_39_DFFSR_3 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_45_DFFSR_87 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_6_DFFSR_232 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_33_DFFSR_159 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_47_DFFSR_263 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_23_DFFSR_162 BUFX2_99/A DFFSR_92/S FILL
XFILL_4_NAND3X1_143 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_37_DFFSR_266 INVX1_67/gnd DFFSR_201/S FILL
XFILL_29_DFFSR_37 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_1_DFFSR_84 BUFX2_99/A DFFSR_7/S FILL
XFILL_1_INVX1_31 INVX1_1/gnd DFFSR_53/S FILL
XFILL_18_DFFSR_77 BUFX2_98/A DFFSR_32/S FILL
XFILL_8_NAND3X1_6 BUFX2_99/A DFFSR_92/S FILL
XFILL_24_DFFPOSX1_3 INVX1_39/gnd DFFSR_34/S FILL
XFILL_13_DFFSR_165 BUFX2_72/gnd DFFSR_201/S FILL
XOAI21X1_101 DFFSR_208/S INVX1_199/Y NAND2X1_132/Y XOR2X1_1/gnd DFFSR_273/D DFFSR_208/S
+ OAI21X1
XFILL_27_DFFSR_269 INVX1_67/gnd DFFSR_201/S FILL
XFILL_23_DFFPOSX1_6 AND2X2_38/B DFFSR_23/S FILL
XFILL_9_DFFPOSX1_17 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_6_NAND2X1_179 INVX1_1/gnd DFFSR_97/S FILL
XFILL_17_DFFSR_272 INVX1_3/gnd DFFSR_23/S FILL
XFILL_22_DFFPOSX1_9 INVX1_67/gnd DFFSR_201/S FILL
XFILL_0_BUFX2_22 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_9_DFFSR_159 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_18_DFFPOSX1_36 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_10_NOR3X1_1 INVX1_3/gnd DFFSR_79/S FILL
XFILL_50_DFFSR_190 INVX1_39/gnd DFFSR_34/S FILL
XFILL_34_1_1 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_40_DFFSR_193 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_2_INVX1_136 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_9_DFFSR_91 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_37_DFFSR_44 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_26_DFFSR_84 BUFX2_99/A DFFSR_7/S FILL
XFILL_3_DFFSR_269 INVX1_67/gnd DFFSR_201/S FILL
XFILL_2_NAND3X1_239 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_30_DFFSR_196 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_32_3_2 INVX1_1/gnd DFFSR_97/S FILL
XFILL_20_DFFSR_199 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_10_DFFSR_34 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_10_DFFSR_202 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_3_NAND3X1_173 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_5_NOR2X1_78 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_43_DFFSR_120 INVX1_3/gnd DFFSR_23/S FILL
XFILL_8_DFFPOSX1_47 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_34_DFFSR_91 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_45_DFFSR_51 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_6_DFFSR_196 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_12_XNOR2X1_2 BUFX2_98/A DFFSR_6/S FILL
XFILL_33_DFFSR_123 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_47_DFFSR_227 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_23_DFFSR_126 BUFX2_99/A DFFSR_7/S FILL
XFILL_4_NAND3X1_107 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_37_DFFSR_230 INVX1_67/gnd DFFSR_201/S FILL
XFILL_1_DFFSR_48 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_2_AND2X2_40 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_18_DFFSR_41 BUFX2_98/A DFFSR_6/S FILL
XFILL_13_DFFSR_129 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_5_BUFX2_76 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_27_DFFSR_233 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_6_NAND2X1_143 INVX1_67/gnd DFFSR_201/S FILL
XFILL_3_AOI21X1_8 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_17_DFFSR_236 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_6_DFFSR_6 BUFX2_79/A DFFSR_6/S FILL
XFILL_42_DFFSR_98 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_9_DFFSR_123 XOR2X1_4/gnd DFFSR_97/S FILL
XNAND2X1_179 NOR2X1_81/Y XOR2X1_14/Y INVX1_1/gnd NAND2X1_179/Y DFFSR_97/S NAND2X1
XFILL_50_DFFSR_154 BUFX2_99/A DFFSR_7/S FILL
XFILL_8_AOI21X1_71 BUFX2_99/A DFFSR_92/S FILL
XFILL_3_AND2X2_7 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_2_INVX1_100 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_40_DFFSR_157 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_9_DFFSR_55 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_26_DFFSR_48 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_15_DFFSR_88 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_3_DFFSR_233 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_2_NAND3X1_203 INVX1_1/gnd DFFSR_97/S FILL
XFILL_30_DFFSR_160 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_44_DFFSR_264 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_20_DFFSR_163 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_4_OR2X2_6 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_34_DFFSR_267 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_5_NAND3X1_7 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_10_DFFSR_166 AND2X2_38/B DFFSR_59/S FILL
XFILL_24_DFFSR_270 INVX1_39/gnd DFFSR_54/S FILL
XFILL_3_NAND3X1_137 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_5_NOR2X1_42 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_14_DFFSR_273 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_8_DFFPOSX1_11 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_45_DFFSR_15 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_34_DFFSR_55 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_5_NAND2X1_173 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_23_DFFSR_95 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_6_DFFSR_160 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_12_DFFPOSX1_3 INVX1_39/gnd DFFSR_34/S FILL
XFILL_47_DFFSR_191 INVX1_67/gnd DFFSR_175/S FILL
XFILL_11_DFFPOSX1_6 AND2X2_38/B DFFSR_23/S FILL
XFILL_1_DFFSR_12 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_37_DFFSR_194 DFFSR_1/gnd DFFSR_81/S FILL
XBUFX2_80 BUFX2_98/A BUFX2_79/A BUFX2_80/Y DFFSR_6/S BUFX2
XFILL_10_DFFPOSX1_9 INVX1_67/gnd DFFSR_201/S FILL
XFILL_17_DFFPOSX1_30 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_5_BUFX2_40 INVX1_1/gnd DFFSR_97/S FILL
XFILL_0_DFFSR_270 INVX1_39/gnd DFFSR_54/S FILL
XFILL_27_DFFSR_197 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_6_NAND2X1_107 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_17_DFFSR_200 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_1_NAND3X1_233 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_51_DFFSR_6 BUFX2_79/A DFFSR_6/S FILL
XFILL_3_INVX1_96 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_42_DFFSR_62 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_9_AOI21X1_32 DFFSR_62/gnd DFFSR_208/S FILL
XNAND2X1_143 NAND2X1_143/A DFFSR_175/S INVX1_67/gnd AOI21X1_47/B DFFSR_201/S NAND2X1
XFILL_2_NOR2X1_79 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_50_DFFSR_118 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_8_AOI21X1_35 INVX1_39/gnd DFFSR_54/S FILL
XFILL_27_DFFPOSX1_19 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_40_DFFSR_121 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_9_DFFSR_19 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_7_AOI21X1_38 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_26_DFFSR_12 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_15_DFFSR_52 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_3_DFFSR_197 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_2_NAND3X1_167 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_2_BUFX2_87 INVX1_1/gnd DFFSR_53/S FILL
XFILL_30_DFFSR_124 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_6_AOI21X1_41 INVX1_39/gnd DFFSR_34/S FILL
XFILL_44_DFFSR_228 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_9_AND2X2_38 AND2X2_38/B DFFSR_59/S FILL
XFILL_7_DFFPOSX1_41 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_20_DFFSR_127 BUFX2_99/A DFFSR_92/S FILL
XFILL_5_AOI21X1_44 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_34_DFFSR_231 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_10_DFFSR_130 BUFX2_79/A DFFSR_6/S FILL
XAOI21X1_41 OAI21X1_74/Y AOI21X1_41/B AOI21X1_40/Y INVX1_39/gnd AND2X2_40/A DFFSR_34/S
+ AOI21X1
XFILL_4_AOI21X1_47 INVX1_67/gnd DFFSR_175/S FILL
XFILL_24_DFFSR_234 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_50_DFFSR_69 BUFX2_98/A DFFSR_32/S FILL
XFILL_0_AOI21X1_9 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_3_NAND3X1_101 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_3_AOI21X1_50 INVX1_67/gnd DFFSR_175/S FILL
XFILL_14_DFFSR_237 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_20_3 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_2_AOI21X1_53 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_33_4_0 INVX1_1/gnd DFFSR_53/S FILL
XFILL_34_DFFSR_19 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_6_DFFSR_66 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_5_NAND2X1_137 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_12_DFFSR_99 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_1_AOI21X1_56 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_23_DFFSR_59 AND2X2_38/B DFFSR_59/S FILL
XFILL_6_DFFSR_124 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_47_DFFSR_155 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_31_6_1 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_0_AOI21X1_59 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_37_DFFSR_158 INVX1_3/gnd DFFSR_23/S FILL
XBUFX2_44 INVX1_59/Y INVX1_3/gnd DFFSR_7/R DFFSR_79/S BUFX2
XFILL_0_DFFSR_234 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_27_DFFSR_161 INVX1_67/gnd DFFSR_175/S FILL
XFILL_3_OAI21X1_119 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_41_DFFSR_265 INVX1_67/gnd DFFSR_175/S FILL
XFILL_26_DFFPOSX1_49 BUFX2_99/A DFFSR_92/S FILL
XFILL_3_INVX1_208 INVX1_39/gnd DFFSR_34/S FILL
XFILL_17_DFFSR_164 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_17_DFFSR_4 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_31_DFFSR_268 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_8_OAI21X1_83 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_1_NAND3X1_197 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_2_NAND3X1_8 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_7_OAI21X1_86 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_21_DFFSR_271 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_31_DFFSR_66 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_42_DFFSR_26 BUFX2_79/A DFFSR_6/S FILL
XFILL_3_INVX1_60 INVX1_39/gnd DFFSR_34/S FILL
XNAND2X1_107 NOR2X1_72/Y INVX1_176/Y OR2X2_3/gnd NAND2X1_107/Y DFFSR_60/S NAND2X1
XFILL_2_NOR2X1_43 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_6_OAI21X1_89 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_11_DFFSR_274 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_5_OAI21X1_92 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_1_BUFX2_5 AND2X2_38/B DFFSR_59/S FILL
XFILL_15_DFFSR_16 DFFSR_28/gnd DFFSR_3/S FILL
XOAI21X1_89 DFFSR_60/S INVX1_185/Y OAI21X1_89/C OR2X2_3/gnd DFFSR_261/D DFFSR_60/S
+ OAI21X1
XFILL_3_DFFSR_161 INVX1_67/gnd DFFSR_175/S FILL
XFILL_2_NAND3X1_131 AND2X2_38/B DFFSR_59/S FILL
XFILL_4_OAI21X1_95 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_2_BUFX2_51 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_44_DFFSR_192 INVX1_1/gnd DFFSR_97/S FILL
XFILL_3_OAI21X1_98 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_7_DFFSR_268 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_4_NAND2X1_167 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_34_DFFSR_195 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_4_AOI21X1_11 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_24_DFFSR_198 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_50_DFFSR_33 BUFX2_98/A DFFSR_32/S FILL
XFILL_39_DFFSR_73 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_14_DFFSR_201 INVX1_67/gnd DFFSR_201/S FILL
XFILL_3_AOI21X1_14 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_2_AOI21X1_17 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_16_DFFPOSX1_24 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_6_DFFSR_30 BUFX2_98/A DFFSR_32/S FILL
XFILL_41_1_1 BUFX2_98/A DFFSR_32/S FILL
XFILL_5_NAND2X1_101 INVX1_39/gnd DFFSR_54/S FILL
XFILL_12_DFFSR_63 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_23_DFFSR_23 AND2X2_38/B DFFSR_23/S FILL
XFILL_1_AOI21X1_20 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_0_DFFPOSX1_3 INVX1_39/gnd DFFSR_34/S FILL
XFILL_47_DFFSR_119 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_0_NAND3X1_227 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_0_AOI21X1_23 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_39_3_2 BUFX2_79/A DFFSR_6/S FILL
XFILL_37_DFFSR_122 BUFX2_79/A DFFSR_7/S FILL
XFILL_0_DFFSR_198 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_51_DFFSR_226 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_27_DFFSR_125 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_9_OAI21X1_44 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_3_INVX1_172 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_41_DFFSR_229 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_26_DFFPOSX1_13 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_47_DFFSR_80 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_6_AND2X2_39 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_17_DFFSR_128 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_1_NAND3X1_161 AND2X2_38/B DFFSR_23/S FILL
XFILL_8_OAI21X1_47 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_31_DFFSR_232 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_7_AOI21X1_7 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_21_DFFSR_235 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_7_OAI21X1_50 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_6_NAND2X1_68 AND2X2_38/B DFFSR_23/S FILL
XFILL_20_DFFSR_70 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_3_INVX1_24 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_31_DFFSR_30 BUFX2_98/A DFFSR_32/S FILL
XFILL_3_DFFSR_77 BUFX2_98/A DFFSR_32/S FILL
XFILL_6_DFFPOSX1_35 INVX1_39/gnd DFFSR_54/S FILL
XFILL_5_NAND2X1_71 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_6_OAI21X1_53 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_11_DFFSR_238 BUFX2_72/gnd DFFSR_276/S FILL
XNAND2X1_68 AND2X2_31/Y AND2X2_32/Y AND2X2_38/B OAI21X1_38/C DFFSR_23/S NAND2X1
XFILL_4_NAND2X1_74 AND2X2_38/B DFFSR_59/S FILL
XFILL_5_OAI21X1_56 DFFSR_46/gnd DFFSR_54/S FILL
XOAI21X1_53 OAI21X1_53/A OAI21X1_53/B OAI21X1_53/C XOR2X1_1/gnd OAI21X1_53/Y DFFSR_151/S
+ OAI21X1
XFILL_3_DFFSR_125 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_2_BUFX2_15 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_42_3 BUFX2_98/A DFFSR_32/S FILL
XFILL_3_NAND2X1_77 AND2X2_38/B DFFSR_23/S FILL
XFILL_4_OAI21X1_59 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_7_XOR2X1_7 BUFX2_98/A DFFSR_6/S FILL
XFILL_44_DFFSR_156 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_10_AOI22X1_3 INVX1_1/gnd DFFSR_97/S FILL
XFILL_3_OAI21X1_62 INVX1_3/gnd DFFSR_79/S FILL
XFILL_2_NAND2X1_80 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_7_DFFSR_232 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_4_NAND2X1_131 INVX1_3/gnd DFFSR_79/S FILL
XFILL_34_DFFSR_159 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_2_OAI21X1_65 INVX1_1/gnd DFFSR_53/S FILL
XFILL_1_NAND2X1_83 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_48_DFFSR_263 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_24_DFFSR_162 BUFX2_99/A DFFSR_92/S FILL
XFILL_1_OAI21X1_68 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_0_NAND2X1_86 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_38_DFFSR_266 INVX1_67/gnd DFFSR_201/S FILL
XFILL_39_DFFSR_37 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_0_INVX1_71 BUFX2_79/A DFFSR_6/S FILL
XFILL_0_INVX1_209 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_28_DFFSR_77 BUFX2_98/A DFFSR_32/S FILL
XFILL_14_DFFSR_165 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_9_NAND3X1_6 BUFX2_99/A DFFSR_92/S FILL
XFILL_28_DFFSR_269 INVX1_67/gnd DFFSR_201/S FILL
XFILL_0_OAI21X1_71 INVX1_3/gnd DFFSR_79/S FILL
XFILL_2_OAI21X1_113 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_25_DFFPOSX1_43 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_18_DFFSR_272 INVX1_3/gnd DFFSR_23/S FILL
XFILL_12_DFFSR_27 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_0_NAND3X1_191 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_5_DFFSR_3 OR2X2_4/gnd DFFSR_3/S FILL
XDFFSR_7 DFFSR_7/Q DFFSR_7/CLK DFFSR_7/R DFFSR_7/S DFFSR_7/D BUFX2_79/A DFFSR_7/S
+ DFFSR
XFILL_0_DFFSR_162 BUFX2_99/A DFFSR_92/S FILL
XDFFSR_272 DFFSR_272/Q CLKBUF1_45/Y DFFSR_266/R DFFSR_23/S DFFSR_272/D INVX1_3/gnd
+ DFFSR_23/S DFFSR
XFILL_41_DFFSR_193 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_3_INVX1_136 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_47_DFFSR_44 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_36_DFFSR_84 BUFX2_99/A DFFSR_7/S FILL
XFILL_4_DFFSR_269 INVX1_67/gnd DFFSR_201/S FILL
XFILL_8_OAI21X1_11 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_31_DFFSR_196 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_1_NAND3X1_125 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_6_NAND2X1_32 INVX1_3/gnd DFFSR_79/S FILL
XFILL_7_OAI21X1_14 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_21_DFFSR_199 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_3_DFFSR_41 BUFX2_98/A DFFSR_6/S FILL
XFILL_20_DFFSR_34 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_3_NAND2X1_161 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_5_NAND2X1_35 INVX1_67/gnd DFFSR_201/S FILL
XFILL_6_OAI21X1_17 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_11_DFFSR_202 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_3_OR2X2_3 OR2X2_3/gnd DFFSR_4/S FILL
XNAND2X1_32 AND2X2_18/B NOR2X1_30/Y INVX1_3/gnd OAI22X1_45/B DFFSR_79/S NAND2X1
XFILL_5_OAI21X1_20 AND2X2_38/B DFFSR_23/S FILL
XFILL_4_NAND2X1_38 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_6_NOR2X1_78 NOR3X1_6/gnd DFFSR_91/S FILL
XOAI21X1_17 AOI21X1_1/A AOI21X1_1/B INVX1_119/Y DFFSR_46/gnd AOI21X1_1/C DFFSR_62/S
+ OAI21X1
XFILL_3_NAND2X1_41 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_4_OAI21X1_23 INVX1_67/gnd DFFSR_201/S FILL
XDFFPOSX1_35 NAND2X1_144/A CLKBUF1_49/Y AOI21X1_48/Y INVX1_39/gnd DFFSR_54/S DFFPOSX1
XFILL_44_DFFSR_120 INVX1_3/gnd DFFSR_23/S FILL
XFILL_29_DFFSR_7 BUFX2_79/A DFFSR_7/S FILL
XFILL_13_XOR2X1_4 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_3_OAI21X1_26 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_2_NAND2X1_44 INVX1_39/gnd DFFSR_34/S FILL
XFILL_15_DFFPOSX1_18 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_7_DFFSR_196 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_13_XNOR2X1_2 BUFX2_98/A DFFSR_6/S FILL
XFILL_44_DFFSR_91 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_34_DFFSR_123 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_2_OAI21X1_29 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_1_NAND2X1_47 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_48_DFFSR_227 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_13_1_2 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_24_DFFSR_126 BUFX2_99/A DFFSR_7/S FILL
XFILL_1_OAI21X1_32 AND2X2_38/B DFFSR_59/S FILL
XFILL_0_NAND2X1_50 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_38_DFFSR_230 INVX1_67/gnd DFFSR_201/S FILL
XFILL_0_INVX1_35 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_0_DFFSR_88 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_0_INVX1_173 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_3_AND2X2_40 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_28_DFFSR_41 BUFX2_98/A DFFSR_6/S FILL
XFILL_17_DFFSR_81 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_14_DFFSR_129 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_28_DFFSR_233 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_0_OAI21X1_35 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_4_AOI21X1_8 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_18_DFFSR_236 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_0_NAND3X1_155 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_50_DFFSR_3 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_5_DFFPOSX1_29 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_0_DFFSR_126 BUFX2_99/A DFFSR_7/S FILL
XDFFSR_236 DFFSR_236/Q CLKBUF1_21/Y BUFX2_68/Y DFFSR_62/S DFFSR_228/Q DFFSR_62/gnd
+ DFFSR_62/S DFFSR
XFILL_6_AOI22X1_10 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_3_INVX1_100 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_41_DFFSR_157 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_36_DFFSR_48 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_25_DFFSR_88 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_8_DFFSR_95 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_5_AOI22X1_13 AND2X2_38/B DFFSR_23/S FILL
XFILL_4_DFFSR_233 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_31_DFFSR_160 XOR2X1_4/gnd DFFSR_97/S FILL
XAOI22X1_10 NOR3X1_4/Y DFFSR_234/D DFFSR_218/Q NOR3X1_3/Y NOR3X1_6/gnd NAND3X1_79/C
+ DFFSR_91/S AOI22X1
XFILL_45_DFFSR_264 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_4_AOI22X1_16 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_21_DFFSR_163 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_40_4_0 BUFX2_98/A DFFSR_6/S FILL
XFILL_14_DFFPOSX1_48 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_35_DFFSR_267 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_3_AOI22X1_19 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_3_NAND2X1_125 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_6_NAND3X1_7 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_11_DFFSR_166 AND2X2_38/B DFFSR_59/S FILL
XFILL_25_DFFSR_270 INVX1_39/gnd DFFSR_54/S FILL
XFILL_2_AOI22X1_22 INVX1_3/gnd DFFSR_79/S FILL
XINVX1_9 INVX1_9/A BUFX2_99/A INVX1_9/Y DFFSR_7/S INVX1
XFILL_6_NOR2X1_42 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_38_6_1 BUFX2_79/A DFFSR_7/S FILL
XFILL_1_AOI22X1_25 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_15_DFFSR_273 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_11_OAI22X1_43 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_0_AOI22X1_28 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_10_OAI22X1_46 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_44_DFFSR_55 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_33_DFFSR_95 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_1_OAI21X1_107 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_7_DFFSR_160 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_24_DFFPOSX1_37 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_1_NAND2X1_11 BUFX2_98/A DFFSR_6/S FILL
XFILL_48_DFFSR_191 INVX1_67/gnd DFFSR_175/S FILL
XFILL_8_NAND3X1_67 XOR2X1_1/gnd DFFSR_151/S FILL
XAND2X2_4 OR2X2_1/A OR2X2_1/B XOR2X1_4/gnd AND2X2_4/Y DFFSR_97/S AND2X2
XFILL_9_OAI22X1_49 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_0_NAND2X1_14 BUFX2_98/A DFFSR_32/S FILL
XFILL_0_INVX1_137 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_8_NAND3X1_240 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_0_DFFSR_52 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_38_DFFSR_194 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_17_DFFSR_45 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_7_NAND3X1_70 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_8_OAI22X1_52 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_4_BUFX2_80 BUFX2_79/A DFFSR_6/S FILL
XFILL_1_DFFSR_270 INVX1_39/gnd DFFSR_54/S FILL
XFILL_28_DFFSR_197 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_6_NAND3X1_73 INVX1_1/gnd DFFSR_97/S FILL
XFILL_18_DFFSR_200 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_5_NAND3X1_76 INVX1_1/gnd DFFSR_53/S FILL
XFILL_0_NAND3X1_119 DFFSR_46/gnd DFFSR_54/S FILL
XNAND3X1_73 DFFSR_170/Q BUFX2_30/Y BUFX2_26/Y INVX1_1/gnd NAND3X1_73/Y DFFSR_97/S
+ NAND3X1
XFILL_4_NAND3X1_79 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_16_DFFSR_1 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_3_NOR2X1_79 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_3_NAND3X1_82 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_2_NAND2X1_155 BUFX2_79/A DFFSR_7/S FILL
XDFFSR_200 DFFSR_208/D CLKBUF1_14/Y BUFX2_64/Y DFFSR_62/S DFFSR_200/D DFFSR_62/gnd
+ DFFSR_62/S DFFSR
XFILL_41_DFFSR_121 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_2_NAND3X1_85 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_36_DFFSR_12 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_25_DFFSR_52 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_8_DFFSR_59 AND2X2_38/B DFFSR_59/S FILL
XFILL_14_DFFSR_92 BUFX2_99/A DFFSR_92/S FILL
XFILL_10_XNOR2X1_3 INVX1_1/gnd DFFSR_97/S FILL
XFILL_4_DFFSR_197 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_31_DFFSR_124 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_1_NAND3X1_88 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_0_BUFX2_2 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_45_DFFSR_228 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_21_DFFSR_127 BUFX2_99/A DFFSR_92/S FILL
XFILL_0_NAND3X1_91 AND2X2_38/B DFFSR_59/S FILL
XFILL_14_DFFPOSX1_12 AND2X2_38/B DFFSR_23/S FILL
XFILL_35_DFFSR_231 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_0_AND2X2_41 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_48_1_1 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_11_DFFSR_130 BUFX2_79/A DFFSR_6/S FILL
XFILL_25_DFFSR_234 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_1_AOI21X1_9 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_15_DFFSR_237 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_46_3_2 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_10_OAI22X1_10 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_44_DFFSR_19 DFFSR_28/gnd DFFSR_8/S FILL
XINVX1_93 INVX1_93/A INVX1_3/gnd INVX1_93/Y DFFSR_23/S INVX1
XFILL_22_DFFSR_99 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_33_DFFSR_59 AND2X2_38/B DFFSR_59/S FILL
XFILL_7_DFFSR_124 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_48_DFFSR_155 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_8_NAND3X1_31 BUFX2_79/A DFFSR_6/S FILL
XFILL_9_OAI22X1_13 INVX1_1/gnd DFFSR_53/S FILL
XFILL_0_DFFSR_16 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_8_NAND3X1_204 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_38_DFFSR_158 INVX1_3/gnd DFFSR_23/S FILL
XFILL_0_INVX1_101 OR2X2_1/gnd DFFSR_51/S FILL
XINVX1_211 INVX1_211/A BUFX2_8/gnd NOR2X1_77/A DFFSR_81/S INVX1
XFILL_7_NAND3X1_34 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_1_DFFSR_234 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_4_BUFX2_44 INVX1_3/gnd DFFSR_79/S FILL
XFILL_8_OAI22X1_16 AND2X2_38/B DFFSR_59/S FILL
XFILL_28_DFFSR_161 INVX1_67/gnd DFFSR_175/S FILL
XFILL_4_DFFPOSX1_23 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_42_DFFSR_265 INVX1_67/gnd DFFSR_175/S FILL
XFILL_4_INVX1_208 INVX1_39/gnd DFFSR_34/S FILL
XFILL_7_OAI22X1_19 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_6_NAND3X1_37 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_18_DFFSR_164 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_32_DFFSR_268 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_6_OAI22X1_22 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_5_NAND3X1_40 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_3_NAND3X1_8 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_14_2_0 INVX1_39/gnd DFFSR_54/S FILL
XNAND3X1_37 DFFSR_13/Q BUFX2_20/Y BUFX2_14/Y OR2X2_4/gnd NAND3X1_37/Y DFFSR_32/S NAND3X1
XFILL_4_NAND3X1_43 BUFX2_99/A DFFSR_7/S FILL
XFILL_22_DFFSR_271 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_41_DFFSR_66 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_5_OAI22X1_25 INVX1_39/gnd DFFSR_54/S FILL
XFILL_3_NOR2X1_43 DFFSR_34/gnd DFFSR_34/S FILL
XOAI22X1_22 INVX1_52/Y OAI22X1_7/B INVX1_53/Y OAI22X1_7/D DFFSR_8/gnd NOR2X1_27/B
+ DFFSR_60/S OAI22X1
XFILL_13_DFFPOSX1_42 INVX1_39/gnd DFFSR_34/S FILL
XFILL_12_DFFSR_274 BUFX2_72/gnd DFFSR_276/S FILL
XDFFSR_164 DFFSR_164/Q CLKBUF1_21/Y BUFX2_60/Y DFFSR_216/S INVX1_87/A OR2X2_2/gnd
+ DFFSR_216/S DFFSR
XFILL_3_NAND3X1_46 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_4_OAI22X1_28 INVX1_3/gnd DFFSR_23/S FILL
XFILL_2_NAND2X1_119 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_12_4_1 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_2_NAND3X1_49 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_3_OAI22X1_31 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_25_DFFSR_16 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_8_DFFSR_23 AND2X2_38/B DFFSR_23/S FILL
XFILL_4_DFFSR_161 INVX1_67/gnd DFFSR_175/S FILL
XFILL_14_DFFSR_56 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_1_BUFX2_91 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_1_NAND3X1_52 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_2_OAI22X1_34 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_45_DFFSR_192 INVX1_1/gnd DFFSR_97/S FILL
XFILL_10_6_2 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_0_NAND3X1_55 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_1_OAI22X1_37 INVX1_3/gnd DFFSR_23/S FILL
XFILL_8_DFFSR_268 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_35_DFFSR_195 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_0_OAI21X1_101 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_23_DFFPOSX1_31 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_0_OAI22X1_40 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_25_DFFSR_198 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_49_DFFSR_73 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_7_4 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_15_DFFSR_201 INVX1_67/gnd DFFSR_201/S FILL
XFILL_7_NAND3X1_234 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_5_DFFSR_70 DFFSR_28/gnd DFFSR_8/S FILL
XINVX1_57 DFFSR_24/D BUFX2_98/A INVX1_57/Y DFFSR_32/S INVX1
XFILL_22_DFFSR_63 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_33_DFFSR_23 AND2X2_38/B DFFSR_23/S FILL
XFILL_0_NOR2X1_80 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_48_DFFSR_119 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_38_DFFSR_122 BUFX2_79/A DFFSR_7/S FILL
XINVX1_175 INVX1_175/A BUFX2_99/A INVX1_175/Y DFFSR_7/S INVX1
XFILL_8_NAND3X1_168 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_1_DFFSR_198 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_28_DFFSR_125 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_1_NAND2X1_149 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_4_INVX1_172 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_42_DFFSR_229 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_7_AND2X2_39 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_18_DFFSR_128 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_32_DFFSR_232 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_8_AOI21X1_7 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_22_DFFSR_235 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_9_NAND3X1_102 INVX1_3/gnd DFFSR_23/S FILL
XFILL_30_DFFSR_70 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_41_DFFSR_30 BUFX2_98/A DFFSR_32/S FILL
XFILL_2_INVX1_64 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_12_DFFSR_238 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_3_NAND3X1_10 BUFX2_79/A DFFSR_6/S FILL
XDFFSR_128 BUFX2_89/A DFFSR_83/CLK DFFSR_73/R DFFSR_91/S INVX1_58/A NOR3X1_6/gnd DFFSR_91/S
+ DFFSR
XFILL_2_NAND3X1_13 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_20_1_2 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_14_DFFSR_20 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_4_DFFSR_125 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_1_NAND3X1_16 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_1_BUFX2_55 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_2_0_1 INVX1_67/gnd DFFSR_201/S FILL
XFILL_45_DFFSR_156 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_11_AOI22X1_3 INVX1_1/gnd DFFSR_97/S FILL
XFILL_0_NAND3X1_19 BUFX2_99/A DFFSR_92/S FILL
XFILL_8_DFFSR_232 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_35_DFFSR_159 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_5_NOR3X1_1 INVX1_3/gnd DFFSR_79/S FILL
XFILL_49_DFFSR_263 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_28_DFFSR_4 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_25_DFFSR_162 BUFX2_99/A DFFSR_92/S FILL
XFILL_0_2_2 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_39_DFFSR_266 INVX1_67/gnd DFFSR_201/S FILL
XFILL_49_DFFSR_37 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_38_DFFSR_77 BUFX2_98/A DFFSR_32/S FILL
XFILL_1_INVX1_209 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_15_DFFSR_165 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_7_NAND3X1_198 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_29_DFFSR_269 INVX1_67/gnd DFFSR_201/S FILL
XFILL_0_NAND3X1_9 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_3_DFFPOSX1_17 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_0_NAND2X1_179 INVX1_1/gnd DFFSR_97/S FILL
XDFFSR_74 INVX1_13/A DFFSR_82/CLK DFFSR_35/R DFFSR_5/S DFFSR_66/Q DFFSR_5/gnd DFFSR_5/S
+ DFFSR
XINVX1_21 INVX1_21/A OR2X2_4/gnd INVX1_21/Y DFFSR_32/S INVX1
XFILL_19_DFFSR_272 INVX1_3/gnd DFFSR_23/S FILL
XFILL_5_DFFSR_34 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_22_DFFSR_27 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_11_DFFSR_67 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_0_NOR2X1_44 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_8_NAND3X1_132 AND2X2_38/B DFFSR_23/S FILL
XINVX1_139 INVX1_139/A DFFSR_1/gnd AOI21X1_8/B DFFSR_81/S INVX1
XFILL_47_4_0 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_12_DFFPOSX1_36 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_1_DFFSR_162 BUFX2_99/A DFFSR_92/S FILL
XFILL_42_DFFSR_193 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_1_NAND2X1_113 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_46_DFFSR_84 BUFX2_99/A DFFSR_7/S FILL
XFILL_5_DFFSR_269 INVX1_67/gnd DFFSR_201/S FILL
XFILL_32_DFFSR_196 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_45_6_1 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_22_DFFSR_199 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_2_INVX1_28 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_2_DFFSR_81 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_30_DFFSR_34 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_19_DFFSR_74 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_12_DFFSR_202 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_22_DFFPOSX1_25 BUFX2_79/A DFFSR_6/S FILL
XFILL_1_BUFX2_19 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_6_NAND3X1_228 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_4_INVX1_2 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_45_DFFSR_120 INVX1_3/gnd DFFSR_23/S FILL
XFILL_8_DFFSR_196 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_14_XNOR2X1_2 BUFX2_98/A DFFSR_6/S FILL
XFILL_2_DFFPOSX1_47 XOR2X1_4/gnd DFFSR_91/S FILL
XNOR3X1_5 NOR3X1_5/A NOR3X1_5/B NOR3X1_5/C BUFX2_7/gnd NOR3X1_5/Y DFFSR_216/S NOR3X1
XFILL_35_DFFSR_123 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_49_DFFSR_227 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_25_DFFSR_126 BUFX2_99/A DFFSR_7/S FILL
XFILL_39_DFFSR_230 INVX1_67/gnd DFFSR_201/S FILL
XFILL_1_INVX1_173 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_4_AND2X2_40 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_38_DFFSR_41 BUFX2_98/A DFFSR_6/S FILL
XFILL_27_DFFSR_81 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_15_DFFSR_129 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_7_NAND3X1_162 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_29_DFFSR_233 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_5_AOI21X1_8 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_0_NAND2X1_143 INVX1_67/gnd DFFSR_201/S FILL
XDFFSR_38 DFFSR_46/D DFFSR_7/CLK DFFSR_2/R DFFSR_6/S DFFSR_38/D BUFX2_98/A DFFSR_6/S
+ DFFSR
XFILL_19_DFFSR_236 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_11_DFFSR_31 BUFX2_79/A DFFSR_6/S FILL
XINVX1_103 DFFSR_246/Q INVX1_39/gnd INVX1_103/Y DFFSR_54/S INVX1
XFILL_1_DFFSR_126 BUFX2_99/A DFFSR_7/S FILL
XFILL_42_DFFSR_157 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_46_DFFSR_48 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_51_5 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_35_DFFSR_88 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_5_DFFSR_233 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_32_DFFSR_160 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_46_DFFSR_264 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_53_3_2 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_22_DFFSR_163 DFFSR_1/gnd DFFSR_1/S FILL
XAOI22X1_1 NOR3X1_2/Y DFFSR_97/Q DFFSR_89/Q NOR3X1_1/Y INVX1_1/gnd AOI22X1_1/Y DFFSR_97/S
+ AOI22X1
XFILL_2_DFFSR_45 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_36_DFFSR_267 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_19_DFFSR_38 BUFX2_98/A DFFSR_6/S FILL
XFILL_7_NAND3X1_7 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_6_BUFX2_73 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_12_DFFSR_166 AND2X2_38/B DFFSR_59/S FILL
XFILL_8_OAI21X1_114 AND2X2_38/B DFFSR_59/S FILL
XFILL_26_DFFSR_270 INVX1_39/gnd DFFSR_54/S FILL
XFILL_16_DFFSR_273 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_20_CLKBUF1_28 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_6_NAND3X1_192 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_12_XOR2X1_8 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_19_CLKBUF1_31 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_2_DFFPOSX1_11 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_43_DFFSR_95 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_8_DFFSR_160 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_18_CLKBUF1_34 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_49_DFFSR_191 INVX1_67/gnd DFFSR_175/S FILL
XNAND3X1_228 OAI21X1_77/Y INVX1_177/A NAND2X1_107/Y OR2X2_3/gnd NAND3X1_228/Y DFFSR_4/S
+ NAND3X1
XFILL_4_AND2X2_4 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_21_2_0 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_1_INVX1_137 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_17_CLKBUF1_37 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_39_DFFSR_194 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_16_DFFSR_85 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_27_DFFSR_45 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_2_DFFSR_270 INVX1_39/gnd DFFSR_54/S FILL
XFILL_7_NAND3X1_126 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_16_CLKBUF1_40 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_29_DFFSR_197 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_11_DFFPOSX1_30 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_0_NAND2X1_107 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_19_4_1 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_15_CLKBUF1_43 AND2X2_38/B DFFSR_23/S FILL
XFILL_19_DFFSR_200 DFFSR_62/gnd DFFSR_62/S FILL
XNOR2X1_82 OR2X2_6/A NOR2X1_82/B XOR2X1_4/gnd NOR2X1_82/Y DFFSR_97/S NOR2X1
XFILL_14_CLKBUF1_46 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_1_3_0 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_13_CLKBUF1_49 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_4_NOR2X1_79 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_40_DFFSR_7 BUFX2_79/A DFFSR_7/S FILL
XFILL_17_6_2 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_21_DFFPOSX1_19 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_42_DFFSR_121 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_46_DFFSR_12 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_7_DFFSR_99 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_35_DFFSR_52 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_24_DFFSR_92 BUFX2_99/A DFFSR_92/S FILL
XFILL_11_XNOR2X1_3 INVX1_1/gnd DFFSR_97/S FILL
XFILL_5_DFFSR_197 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_32_DFFSR_124 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_5_NAND3X1_222 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_46_DFFSR_228 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_22_DFFSR_127 BUFX2_99/A DFFSR_92/S FILL
XFILL_1_DFFPOSX1_41 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_36_DFFSR_231 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_1_AND2X2_41 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_12_DFFSR_130 BUFX2_79/A DFFSR_6/S FILL
XFILL_6_BUFX2_37 INVX1_1/gnd DFFSR_97/S FILL
XFILL_26_DFFSR_234 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_11_2 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_2_AOI21X1_9 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_16_DFFSR_237 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_6_NAND3X1_156 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_32_DFFSR_99 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_4_INVX1_93 INVX1_3/gnd DFFSR_23/S FILL
XFILL_43_DFFSR_59 AND2X2_38/B DFFSR_59/S FILL
XFILL_8_DFFSR_124 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_49_DFFSR_155 OR2X2_1/gnd DFFSR_59/S FILL
XNAND3X1_192 AOI21X1_26/C NAND3X1_192/B NAND3X1_192/C OR2X2_2/gnd AOI21X1_25/A DFFSR_216/S
+ NAND3X1
XFILL_39_DFFSR_158 INVX1_3/gnd DFFSR_23/S FILL
XFILL_1_INVX1_101 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_16_DFFSR_49 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_2_DFFSR_234 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_29_DFFSR_161 INVX1_67/gnd DFFSR_175/S FILL
XFILL_3_BUFX2_84 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_43_DFFSR_265 INVX1_67/gnd DFFSR_175/S FILL
XFILL_20_DFFPOSX1_49 BUFX2_99/A DFFSR_92/S FILL
XFILL_19_DFFSR_164 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_33_DFFSR_268 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_27_1_2 INVX1_3/gnd DFFSR_79/S FILL
XNOR2X1_46 NOR2X1_46/A NOR2X1_46/B DFFSR_34/gnd NOR2X1_46/Y DFFSR_1/S NOR2X1
XFILL_4_NAND3X1_8 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_14_CLKBUF1_10 INVX1_67/gnd DFFSR_201/S FILL
XFILL_23_DFFSR_271 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_51_DFFSR_66 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_13_CLKBUF1_13 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_4_NOR2X1_43 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_9_0_1 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_13_DFFSR_274 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_12_CLKBUF1_16 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_7_OAI21X1_108 INVX1_1/gnd DFFSR_53/S FILL
XFILL_35_DFFSR_16 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_7_DFFSR_63 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_7_2_2 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_24_DFFSR_56 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_13_DFFSR_96 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_11_CLKBUF1_19 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_5_DFFSR_161 INVX1_67/gnd DFFSR_175/S FILL
XFILL_5_NAND3X1_186 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_46_DFFSR_192 INVX1_1/gnd DFFSR_97/S FILL
XFILL_10_CLKBUF1_22 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_9_DFFSR_268 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_36_DFFSR_195 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_26_DFFSR_198 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_9_CLKBUF1_25 INVX1_67/gnd DFFSR_201/S FILL
XFILL_16_DFFSR_201 INVX1_67/gnd DFFSR_201/S FILL
XFILL_8_CLKBUF1_28 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_27_DFFSR_1 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_6_NAND3X1_120 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_7_CLKBUF1_31 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_54_4_0 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_10_DFFPOSX1_24 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_32_DFFSR_63 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_4_INVX1_57 BUFX2_98/A DFFSR_32/S FILL
XFILL_43_DFFSR_23 AND2X2_38/B DFFSR_23/S FILL
XFILL_6_CLKBUF1_34 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_1_NOR2X1_80 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_49_DFFSR_119 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_5_CLKBUF1_37 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_52_6_1 BUFX2_77/gnd DFFSR_98/S FILL
XNAND3X1_156 INVX1_151/Y AOI22X1_21/C NAND2X1_74/Y OR2X2_1/gnd AOI21X1_11/A DFFSR_59/S
+ NAND3X1
XFILL_39_DFFSR_122 BUFX2_79/A DFFSR_7/S FILL
XCLKBUF1_34 BUFX2_5/Y BUFX2_72/gnd CLKBUF1_34/Y DFFSR_201/S CLKBUF1
XFILL_16_DFFSR_13 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_4_CLKBUF1_40 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_2_DFFSR_198 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_29_DFFSR_125 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_3_BUFX2_48 AND2X2_38/B DFFSR_59/S FILL
XFILL_43_DFFSR_229 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_8_AND2X2_39 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_3_CLKBUF1_43 AND2X2_38/B DFFSR_23/S FILL
XFILL_19_DFFSR_128 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_20_DFFPOSX1_13 BUFX2_8/gnd DFFSR_81/S FILL
XXNOR2X1_1 XNOR2X1_1/A XNOR2X1_1/B BUFX2_8/gnd INVX1_164/A DFFSR_51/S XNOR2X1
XFILL_33_DFFSR_232 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_2_CLKBUF1_46 OR2X2_3/gnd DFFSR_4/S FILL
XNOR2X1_10 OAI22X1_6/Y OAI21X1_2/Y BUFX2_98/A NOR2X1_10/Y DFFSR_32/S NOR2X1
XFILL_9_AOI21X1_7 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_23_DFFSR_235 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_1_CLKBUF1_49 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_4_NAND3X1_216 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_51_DFFSR_30 BUFX2_98/A DFFSR_32/S FILL
XFILL_40_DFFSR_70 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_13_DFFSR_238 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_0_DFFPOSX1_35 INVX1_39/gnd DFFSR_54/S FILL
XFILL_33_2 INVX1_1/gnd DFFSR_97/S FILL
XFILL_7_DFFSR_27 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_13_DFFSR_60 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_24_DFFSR_20 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_5_DFFSR_125 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_0_BUFX2_95 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_46_DFFSR_156 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_5_NAND3X1_150 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_9_DFFSR_232 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_36_DFFSR_159 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_6_NOR2X1_8 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_50_DFFSR_263 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_26_DFFSR_162 BUFX2_99/A DFFSR_92/S FILL
XFILL_40_DFFSR_266 INVX1_67/gnd DFFSR_201/S FILL
XFILL_48_DFFSR_77 BUFX2_98/A DFFSR_32/S FILL
XFILL_2_INVX1_209 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_16_DFFSR_165 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_30_DFFSR_269 INVX1_67/gnd DFFSR_201/S FILL
XFILL_1_NAND3X1_9 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_20_DFFSR_272 INVX1_3/gnd DFFSR_23/S FILL
XFILL_32_DFFSR_27 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_4_DFFSR_74 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_4_INVX1_21 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_21_DFFSR_67 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_19_DFFPOSX1_43 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_1_NOR2X1_44 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_10_DFFSR_275 BUFX2_99/A DFFSR_92/S FILL
XNAND3X1_120 NOR2X1_53/Y NOR2X1_54/Y NOR2X1_55/Y BUFX2_8/gnd XOR2X1_15/B DFFSR_51/S
+ NAND3X1
XFILL_3_NAND3X1_246 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_3_BUFX2_12 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_2_DFFSR_162 BUFX2_99/A DFFSR_92/S FILL
XFILL_8_XOR2X1_4 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_43_DFFSR_193 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_6_OAI21X1_102 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_6_DFFSR_269 INVX1_67/gnd DFFSR_201/S FILL
XFILL_33_DFFSR_196 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_2_CLKBUF1_10 INVX1_67/gnd DFFSR_201/S FILL
XFILL_1_CLKBUF1_13 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_4_NAND3X1_180 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_23_DFFSR_199 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_1_INVX1_68 INVX1_67/gnd DFFSR_201/S FILL
XFILL_29_DFFSR_74 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_40_DFFSR_34 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_0_CLKBUF1_16 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_13_DFFSR_202 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_13_DFFSR_24 BUFX2_98/A DFFSR_6/S FILL
XFILL_28_2_0 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_0_BUFX2_59 AND2X2_38/B DFFSR_23/S FILL
XFILL_46_DFFSR_120 INVX1_3/gnd DFFSR_23/S FILL
XFILL_5_NAND3X1_114 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_15_XNOR2X1_2 BUFX2_98/A DFFSR_6/S FILL
XFILL_9_DFFSR_196 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_36_DFFSR_123 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_4_NOR3X1_5 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_50_DFFSR_227 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_26_4_1 INVX1_3/gnd DFFSR_23/S FILL
XFILL_18_DFFSR_8 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_26_DFFSR_126 BUFX2_99/A DFFSR_7/S FILL
XFILL_40_DFFSR_230 INVX1_67/gnd DFFSR_201/S FILL
XFILL_8_3_0 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_2_INVX1_173 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_48_DFFSR_41 BUFX2_98/A DFFSR_6/S FILL
XFILL_37_DFFSR_81 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_5_AND2X2_40 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_16_DFFSR_129 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_30_DFFSR_233 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_24_6_2 AND2X2_38/B DFFSR_59/S FILL
XFILL_6_AOI21X1_8 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_20_DFFSR_236 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_6_5_1 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_4_DFFSR_38 BUFX2_98/A DFFSR_6/S FILL
XFILL_21_DFFSR_31 BUFX2_79/A DFFSR_6/S FILL
XFILL_10_DFFSR_71 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_2_BUFX2_9 AND2X2_38/B DFFSR_59/S FILL
XFILL_10_DFFSR_239 INVX1_39/gnd DFFSR_54/S FILL
XFILL_3_NAND3X1_210 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_2_DFFSR_126 BUFX2_99/A DFFSR_7/S FILL
XFILL_43_DFFSR_157 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_55_2 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_14_XOR2X1_1 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_39_DFFSR_4 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_45_DFFSR_88 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_6_DFFSR_233 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_33_DFFSR_160 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_47_DFFSR_264 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_25_DFFPOSX1_1 INVX1_39/gnd DFFSR_34/S FILL
XFILL_4_NAND3X1_144 AND2X2_38/B DFFSR_59/S FILL
XFILL_23_DFFSR_163 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_1_INVX1_32 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_37_DFFSR_267 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_1_DFFSR_85 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_18_DFFSR_78 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_29_DFFSR_38 BUFX2_98/A DFFSR_6/S FILL
XFILL_24_DFFPOSX1_4 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_8_NAND3X1_7 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_13_DFFSR_166 AND2X2_38/B DFFSR_59/S FILL
XOAI21X1_102 DFFSR_276/S INVX1_200/Y NAND2X1_133/Y BUFX2_72/gnd DFFSR_274/D DFFSR_201/S
+ OAI21X1
XFILL_27_DFFSR_270 INVX1_39/gnd DFFSR_54/S FILL
XFILL_9_DFFPOSX1_18 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_23_DFFPOSX1_7 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_6_NAND2X1_180 INVX1_1/gnd DFFSR_97/S FILL
XFILL_17_DFFSR_273 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_0_BUFX2_23 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_9_DFFSR_160 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_18_DFFPOSX1_37 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_50_DFFSR_191 INVX1_67/gnd DFFSR_175/S FILL
XFILL_10_NOR3X1_2 INVX1_1/gnd DFFSR_53/S FILL
XFILL_34_1_2 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_40_DFFSR_194 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_2_INVX1_137 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_37_DFFSR_45 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_9_DFFSR_92 BUFX2_99/A DFFSR_92/S FILL
XFILL_26_DFFSR_85 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_2_NAND3X1_240 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_3_DFFSR_270 INVX1_39/gnd DFFSR_54/S FILL
XFILL_30_DFFSR_197 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_20_DFFSR_200 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_10_DFFSR_35 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_10_DFFSR_203 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_3_NAND3X1_174 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_5_NOR2X1_79 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_43_DFFSR_121 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_8_DFFPOSX1_48 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_45_DFFSR_52 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_34_DFFSR_92 BUFX2_99/A DFFSR_92/S FILL
XFILL_12_XNOR2X1_3 INVX1_1/gnd DFFSR_97/S FILL
XFILL_6_DFFSR_197 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_33_DFFSR_124 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_47_DFFSR_228 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_23_DFFSR_127 BUFX2_99/A DFFSR_92/S FILL
XFILL_4_NAND3X1_108 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_37_DFFSR_231 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_18_DFFSR_42 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_1_DFFSR_49 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_2_AND2X2_41 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_5_BUFX2_77 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_13_DFFSR_130 BUFX2_79/A DFFSR_6/S FILL
XFILL_27_DFFSR_234 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_3_AOI21X1_9 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_6_NAND2X1_144 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_17_DFFSR_237 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_6_DFFSR_7 BUFX2_79/A DFFSR_7/S FILL
XFILL_42_DFFSR_99 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_9_DFFSR_124 OR2X2_1/gnd DFFSR_59/S FILL
XNAND2X1_180 NAND2X1_180/A NAND2X1_179/Y INVX1_1/gnd OR2X2_6/B DFFSR_97/S NAND2X1
XFILL_50_DFFSR_155 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_3_AND2X2_8 BUFX2_99/A DFFSR_7/S FILL
XFILL_40_DFFSR_158 INVX1_3/gnd DFFSR_23/S FILL
XFILL_9_DFFSR_56 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_2_INVX1_101 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_26_DFFSR_49 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_2_NAND3X1_204 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_15_DFFSR_89 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_3_DFFSR_234 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_30_DFFSR_161 INVX1_67/gnd DFFSR_175/S FILL
XFILL_44_DFFSR_265 INVX1_67/gnd DFFSR_175/S FILL
XFILL_20_DFFSR_164 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_34_DFFSR_268 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_5_NAND3X1_8 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_10_DFFSR_167 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_24_DFFSR_271 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_3_NAND3X1_138 INVX1_67/gnd DFFSR_201/S FILL
XFILL_5_NOR2X1_43 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_14_DFFSR_274 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_8_DFFPOSX1_12 AND2X2_38/B DFFSR_23/S FILL
XFILL_13_DFFPOSX1_1 INVX1_39/gnd DFFSR_34/S FILL
XFILL_5_NAND2X1_174 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_45_DFFSR_16 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_34_DFFSR_56 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_23_DFFSR_96 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_6_DFFSR_161 INVX1_67/gnd DFFSR_175/S FILL
XFILL_12_DFFPOSX1_4 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_47_DFFSR_192 INVX1_1/gnd DFFSR_97/S FILL
XFILL_11_DFFPOSX1_7 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_1_DFFSR_13 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_37_DFFSR_195 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_5_BUFX2_41 BUFX2_77/gnd DFFSR_5/S FILL
XBUFX2_81 BUFX2_79/A BUFX2_79/A BUFX2_81/Y DFFSR_7/S BUFX2
XFILL_0_DFFSR_271 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_17_DFFPOSX1_31 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_27_DFFSR_198 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_6_NAND2X1_108 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_17_DFFSR_201 INVX1_67/gnd DFFSR_201/S FILL
XFILL_1_NAND3X1_234 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_42_DFFSR_63 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_3_INVX1_97 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_2_NOR2X1_80 NOR3X1_6/gnd DFFSR_91/S FILL
XNAND2X1_144 NAND2X1_144/A INVX1_208/Y DFFSR_46/gnd AOI21X1_48/A DFFSR_62/S NAND2X1
XFILL_50_DFFSR_119 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_8_AOI21X1_36 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_27_DFFPOSX1_20 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_40_DFFSR_122 BUFX2_79/A DFFSR_7/S FILL
XFILL_7_AOI21X1_39 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_9_DFFSR_20 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_26_DFFSR_13 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_15_DFFSR_53 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_2_NAND3X1_168 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_3_DFFSR_198 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_30_DFFSR_125 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_2_BUFX2_88 INVX1_3/gnd DFFSR_23/S FILL
XFILL_44_DFFSR_229 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_6_AOI21X1_42 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_20_DFFSR_128 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_7_DFFPOSX1_42 INVX1_39/gnd DFFSR_34/S FILL
XFILL_5_AOI21X1_45 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_34_DFFSR_232 DFFSR_46/gnd DFFSR_54/S FILL
XAOI21X1_42 NAND2X1_99/A NAND2X1_99/B INVX1_169/A DFFSR_34/gnd AOI21X1_42/Y DFFSR_34/S
+ AOI21X1
XFILL_10_DFFSR_131 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_35_2_0 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_4_AOI21X1_48 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_24_DFFSR_235 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_50_DFFSR_70 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_3_NAND3X1_102 INVX1_3/gnd DFFSR_23/S FILL
XFILL_3_AOI21X1_51 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_14_DFFSR_238 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_20_4 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_33_4_1 INVX1_1/gnd DFFSR_53/S FILL
XFILL_2_AOI21X1_54 AND2X2_38/B DFFSR_59/S FILL
XFILL_5_NAND2X1_138 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_23_DFFSR_60 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_34_DFFSR_20 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_6_DFFSR_67 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_1_AOI21X1_57 INVX1_67/gnd DFFSR_201/S FILL
XFILL_6_DFFSR_125 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_47_DFFSR_156 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_0_AOI21X1_60 BUFX2_79/A DFFSR_7/S FILL
XFILL_31_6_2 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_37_DFFSR_159 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_0_DFFSR_235 OR2X2_2/gnd DFFSR_216/S FILL
XBUFX2_45 INVX1_59/Y BUFX2_77/gnd DFFSR_15/R DFFSR_5/S BUFX2
XFILL_27_DFFSR_162 BUFX2_99/A DFFSR_92/S FILL
XFILL_41_DFFSR_266 INVX1_67/gnd DFFSR_201/S FILL
XFILL_9_OAI21X1_81 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_26_DFFPOSX1_50 INVX1_1/gnd DFFSR_53/S FILL
XFILL_3_INVX1_209 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_17_DFFSR_165 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_17_DFFSR_5 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_8_OAI21X1_84 BUFX2_98/A DFFSR_6/S FILL
XFILL_31_DFFSR_269 INVX1_67/gnd DFFSR_201/S FILL
XFILL_1_NAND3X1_198 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_2_NAND3X1_9 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_7_OAI21X1_87 BUFX2_79/A DFFSR_7/S FILL
XFILL_21_DFFSR_272 INVX1_3/gnd DFFSR_23/S FILL
XFILL_42_DFFSR_27 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_3_INVX1_61 INVX1_39/gnd DFFSR_54/S FILL
XFILL_31_DFFSR_67 DFFSR_34/gnd DFFSR_34/S FILL
XNAND2X1_108 NOR2X1_72/Y XNOR2X1_2/Y DFFSR_8/gnd NAND2X1_108/Y DFFSR_60/S NAND2X1
XFILL_2_NOR2X1_44 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_6_OAI21X1_90 BUFX2_98/A DFFSR_32/S FILL
XFILL_11_DFFSR_275 BUFX2_99/A DFFSR_92/S FILL
XFILL_5_OAI21X1_93 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_1_BUFX2_6 BUFX2_79/A DFFSR_6/S FILL
XFILL_15_DFFSR_17 DFFSR_28/gnd DFFSR_3/S FILL
XOAI21X1_90 DFFSR_32/S INVX1_186/Y OAI21X1_90/C BUFX2_98/A DFFSR_262/D DFFSR_32/S
+ OAI21X1
XFILL_2_NAND3X1_132 AND2X2_38/B DFFSR_23/S FILL
XFILL_3_DFFSR_162 BUFX2_99/A DFFSR_92/S FILL
XFILL_4_OAI21X1_96 AND2X2_38/B DFFSR_59/S FILL
XFILL_2_BUFX2_52 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_44_DFFSR_193 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_3_OAI21X1_99 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_7_DFFSR_269 INVX1_67/gnd DFFSR_201/S FILL
XFILL_34_DFFSR_196 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_4_NAND2X1_168 BUFX2_79/A DFFSR_6/S FILL
XFILL_38_DFFSR_1 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_4_AOI21X1_12 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_24_DFFSR_199 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_39_DFFSR_74 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_50_DFFSR_34 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_3_AOI21X1_15 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_14_DFFSR_202 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_1_DFFPOSX1_1 INVX1_39/gnd DFFSR_34/S FILL
XFILL_2_AOI21X1_18 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_16_DFFPOSX1_25 BUFX2_79/A DFFSR_6/S FILL
XFILL_5_NAND2X1_102 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_12_DFFSR_64 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_41_1_2 BUFX2_98/A DFFSR_32/S FILL
XFILL_23_DFFSR_24 BUFX2_98/A DFFSR_6/S FILL
XFILL_6_DFFSR_31 BUFX2_79/A DFFSR_6/S FILL
XFILL_1_AOI21X1_21 INVX1_39/gnd DFFSR_54/S FILL
XFILL_0_DFFPOSX1_4 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_0_NAND3X1_228 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_47_DFFSR_120 INVX1_3/gnd DFFSR_23/S FILL
XFILL_0_AOI21X1_24 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_37_DFFSR_123 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_0_DFFSR_199 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_27_DFFSR_126 BUFX2_99/A DFFSR_7/S FILL
XFILL_41_DFFSR_230 INVX1_67/gnd DFFSR_201/S FILL
XFILL_26_DFFPOSX1_14 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_3_INVX1_173 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_47_DFFSR_81 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_6_AND2X2_40 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_17_DFFSR_129 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_8_OAI21X1_48 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_31_DFFSR_233 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_1_NAND3X1_162 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_7_AOI21X1_8 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_6_NAND2X1_69 INVX1_3/gnd DFFSR_23/S FILL
XFILL_7_OAI21X1_51 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_21_DFFSR_236 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_3_INVX1_25 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_3_DFFSR_78 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_31_DFFSR_31 BUFX2_79/A DFFSR_6/S FILL
XFILL_20_DFFSR_71 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_6_DFFPOSX1_36 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_5_NAND2X1_72 AND2X2_38/B DFFSR_59/S FILL
XFILL_11_DFFSR_239 INVX1_39/gnd DFFSR_54/S FILL
XFILL_6_OAI21X1_54 XOR2X1_1/gnd DFFSR_208/S FILL
XNAND2X1_69 BUFX2_59/Y AND2X2_34/B INVX1_3/gnd OAI21X1_31/C DFFSR_23/S NAND2X1
XFILL_4_NAND2X1_75 INVX1_3/gnd DFFSR_79/S FILL
XFILL_5_OAI21X1_57 DFFSR_34/gnd DFFSR_34/S FILL
XOAI21X1_54 OAI21X1_54/A OAI21X1_54/B OAI21X1_54/C XOR2X1_1/gnd OAI21X1_54/Y DFFSR_208/S
+ OAI21X1
XFILL_42_4 BUFX2_98/A DFFSR_32/S FILL
XFILL_3_DFFSR_126 BUFX2_99/A DFFSR_7/S FILL
XFILL_3_NAND2X1_78 AND2X2_38/B DFFSR_23/S FILL
XFILL_4_OAI21X1_60 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_2_BUFX2_16 BUFX2_98/A DFFSR_32/S FILL
XFILL_7_XOR2X1_8 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_44_DFFSR_157 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_10_AOI22X1_4 BUFX2_99/A DFFSR_92/S FILL
XFILL_2_NAND2X1_81 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_3_OAI21X1_63 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_7_DFFSR_233 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_4_NAND2X1_132 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_34_DFFSR_160 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_48_DFFSR_264 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_2_OAI21X1_66 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_1_NAND2X1_84 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_24_DFFSR_163 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_0_NAND2X1_87 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_1_OAI21X1_69 INVX1_3/gnd DFFSR_23/S FILL
XFILL_28_DFFSR_78 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_39_DFFSR_38 BUFX2_98/A DFFSR_6/S FILL
XFILL_0_INVX1_210 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_0_INVX1_72 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_38_DFFSR_267 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_14_DFFSR_166 AND2X2_38/B DFFSR_59/S FILL
XFILL_0_OAI21X1_72 INVX1_3/gnd DFFSR_23/S FILL
XFILL_28_DFFSR_270 INVX1_39/gnd DFFSR_54/S FILL
XFILL_2_OAI21X1_114 AND2X2_38/B DFFSR_59/S FILL
XFILL_25_DFFPOSX1_44 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_18_DFFSR_273 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_12_DFFSR_28 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_0_NAND3X1_192 OR2X2_2/gnd DFFSR_216/S FILL
XDFFSR_8 DFFSR_8/Q DFFSR_8/CLK DFFSR_8/R DFFSR_8/S DFFSR_8/D DFFSR_8/gnd DFFSR_8/S
+ DFFSR
XFILL_5_DFFSR_4 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_51_DFFSR_191 INVX1_67/gnd DFFSR_175/S FILL
XFILL_0_DFFSR_163 DFFSR_1/gnd DFFSR_1/S FILL
XDFFSR_273 BUFX2_71/A CLKBUF1_15/Y DFFSR_274/R DFFSR_208/S DFFSR_273/D DFFSR_62/gnd
+ DFFSR_208/S DFFSR
XFILL_41_DFFSR_194 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_3_INVX1_137 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_47_DFFSR_45 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_36_DFFSR_85 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_4_DFFSR_270 INVX1_39/gnd DFFSR_54/S FILL
XFILL_8_OAI21X1_12 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_31_DFFSR_197 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_1_NAND3X1_126 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_6_NAND2X1_33 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_7_OAI21X1_15 INVX1_3/gnd DFFSR_79/S FILL
XFILL_21_DFFSR_200 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_3_DFFSR_42 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_20_DFFSR_35 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_3_NAND2X1_162 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_5_NAND2X1_36 INVX1_3/gnd DFFSR_79/S FILL
XFILL_6_OAI21X1_18 INVX1_39/gnd DFFSR_34/S FILL
XFILL_11_DFFSR_203 DFFSR_46/gnd DFFSR_54/S FILL
XNAND2X1_33 NOR3X1_4/B INVX1_63/Y XOR2X1_4/gnd NOR2X1_34/B DFFSR_91/S NAND2X1
XFILL_3_OR2X2_4 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_4_NAND2X1_39 BUFX2_98/A DFFSR_6/S FILL
XFILL_5_OAI21X1_21 AND2X2_38/B DFFSR_59/S FILL
XFILL_6_NOR2X1_79 DFFSR_46/gnd DFFSR_54/S FILL
XOAI21X1_18 AOI21X1_3/B AND2X2_27/B AOI21X1_3/Y INVX1_39/gnd DFFPOSX1_1/D DFFSR_34/S
+ OAI21X1
XFILL_4_OAI21X1_24 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_3_NAND2X1_42 DFFSR_34/gnd DFFSR_34/S FILL
XDFFPOSX1_36 NAND2X1_143/A CLKBUF1_43/Y AOI21X1_46/Y OR2X2_2/gnd DFFSR_175/S DFFPOSX1
XFILL_13_XOR2X1_5 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_44_DFFSR_121 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_3_OAI21X1_27 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_29_DFFSR_8 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_15_DFFPOSX1_19 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_2_NAND2X1_45 INVX1_39/gnd DFFSR_34/S FILL
XFILL_44_DFFSR_92 BUFX2_99/A DFFSR_92/S FILL
XFILL_13_XNOR2X1_3 INVX1_1/gnd DFFSR_97/S FILL
XFILL_7_DFFSR_197 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_34_DFFSR_124 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_1_NAND2X1_48 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_2_OAI21X1_30 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_48_DFFSR_228 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_24_DFFSR_127 BUFX2_99/A DFFSR_92/S FILL
XFILL_5_AND2X2_1 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_0_NAND2X1_51 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_1_OAI21X1_33 INVX1_3/gnd DFFSR_79/S FILL
XFILL_0_INVX1_174 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_0_INVX1_36 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_28_DFFSR_42 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_0_DFFSR_89 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_38_DFFSR_231 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_17_DFFSR_82 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_3_AND2X2_41 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_14_DFFSR_130 BUFX2_79/A DFFSR_6/S FILL
XFILL_0_OAI21X1_36 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_28_DFFSR_234 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_4_AOI21X1_9 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_18_DFFSR_237 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_0_NAND3X1_156 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_9_NAND3X1_211 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_50_DFFSR_4 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_5_DFFPOSX1_30 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_51_DFFSR_155 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_0_DFFSR_127 BUFX2_99/A DFFSR_92/S FILL
XDFFSR_237 DFFSR_245/D CLKBUF1_6/Y BUFX2_66/Y DFFSR_1/S DFFSR_237/D DFFSR_1/gnd DFFSR_1/S
+ DFFSR
XFILL_6_AOI22X1_11 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_41_DFFSR_158 INVX1_3/gnd DFFSR_23/S FILL
XFILL_8_DFFSR_96 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_42_2_0 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_3_INVX1_101 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_36_DFFSR_49 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_25_DFFSR_89 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_5_AOI22X1_14 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_4_DFFSR_234 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_31_DFFSR_161 INVX1_67/gnd DFFSR_175/S FILL
XFILL_45_DFFSR_265 INVX1_67/gnd DFFSR_175/S FILL
XAOI22X1_11 NOR3X1_4/Y DFFSR_235/D DFFSR_219/Q NOR3X1_3/Y BUFX2_7/gnd AOI22X1_11/Y
+ DFFSR_151/S AOI22X1
XFILL_4_AOI22X1_17 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_21_DFFSR_164 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_40_4_1 BUFX2_98/A DFFSR_6/S FILL
XFILL_14_DFFPOSX1_49 BUFX2_99/A DFFSR_92/S FILL
XFILL_35_DFFSR_268 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_6_NAND3X1_8 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_3_AOI22X1_20 INVX1_39/gnd DFFSR_34/S FILL
XFILL_3_NAND2X1_126 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_11_DFFSR_167 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_25_DFFSR_271 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_2_AOI22X1_23 INVX1_39/gnd DFFSR_34/S FILL
XFILL_6_NOR2X1_43 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_15_DFFSR_274 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_38_6_2 BUFX2_79/A DFFSR_7/S FILL
XFILL_1_AOI22X1_26 INVX1_1/gnd DFFSR_97/S FILL
XFILL_11_OAI22X1_44 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_0_AOI22X1_29 INVX1_1/gnd DFFSR_53/S FILL
XFILL_10_OAI22X1_47 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_44_DFFSR_56 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_33_DFFSR_96 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_1_OAI21X1_108 INVX1_1/gnd DFFSR_53/S FILL
XFILL_7_DFFSR_161 INVX1_67/gnd DFFSR_175/S FILL
XFILL_24_DFFPOSX1_38 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_9_NAND3X1_65 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_48_DFFSR_192 INVX1_1/gnd DFFSR_97/S FILL
XFILL_1_NAND2X1_12 INVX1_3/gnd DFFSR_79/S FILL
XFILL_8_NAND3X1_68 BUFX2_7/gnd DFFSR_216/S FILL
XAND2X2_5 BUFX2_19/Y NOR2X1_4/Y DFFSR_8/gnd AND2X2_5/Y DFFSR_8/S AND2X2
XFILL_9_OAI22X1_50 INVX1_3/gnd DFFSR_23/S FILL
XFILL_0_NAND2X1_15 BUFX2_99/A DFFSR_92/S FILL
XFILL_8_NAND3X1_241 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_0_DFFSR_53 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_0_INVX1_138 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_38_DFFSR_195 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_17_DFFSR_46 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_7_NAND3X1_71 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_1_DFFSR_271 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_4_BUFX2_81 BUFX2_79/A DFFSR_7/S FILL
XFILL_28_DFFSR_198 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_6_NAND3X1_74 INVX1_1/gnd DFFSR_97/S FILL
XFILL_18_DFFSR_201 INVX1_67/gnd DFFSR_201/S FILL
XFILL_5_NAND3X1_77 DFFSR_5/gnd DFFSR_5/S FILL
XNAND3X1_74 DFFSR_154/D AND2X2_18/B BUFX2_30/Y INVX1_1/gnd AND2X2_20/B DFFSR_97/S
+ NAND3X1
XFILL_0_NAND3X1_120 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_4_NAND3X1_80 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_16_DFFSR_2 BUFX2_79/A DFFSR_7/S FILL
XFILL_3_NOR2X1_80 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_3_NAND3X1_83 XOR2X1_1/gnd DFFSR_151/S FILL
XDFFSR_201 INVX1_65/A CLKBUF1_34/Y BUFX2_62/Y DFFSR_201/S DFFSR_201/D INVX1_67/gnd
+ DFFSR_201/S DFFSR
XFILL_2_NAND2X1_156 AND2X2_38/B DFFSR_59/S FILL
XFILL_41_DFFSR_122 BUFX2_79/A DFFSR_7/S FILL
XFILL_8_DFFSR_60 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_2_NAND3X1_86 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_14_DFFSR_93 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_36_DFFSR_13 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_25_DFFSR_53 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_4_DFFSR_198 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_10_XNOR2X1_4 BUFX2_98/A DFFSR_6/S FILL
XFILL_31_DFFSR_125 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_1_NAND3X1_89 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_45_DFFSR_229 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_0_BUFX2_3 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_21_DFFSR_128 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_0_NAND3X1_92 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_14_DFFPOSX1_13 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_35_DFFSR_232 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_0_AND2X2_42 INVX1_3/gnd DFFSR_23/S FILL
XFILL_48_1_2 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_11_DFFSR_131 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_25_DFFSR_235 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_24_1 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_15_DFFSR_238 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_10_OAI22X1_11 BUFX2_99/A DFFSR_92/S FILL
XINVX1_94 INVX1_94/A INVX1_67/gnd INVX1_94/Y DFFSR_201/S INVX1
XFILL_33_DFFSR_60 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_44_DFFSR_20 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_7_DFFSR_125 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_9_NAND3X1_29 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_48_DFFSR_156 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_9_OAI22X1_14 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_8_NAND3X1_32 BUFX2_79/A DFFSR_7/S FILL
XFILL_38_DFFSR_159 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_0_DFFSR_17 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_17_DFFSR_10 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_8_NAND3X1_205 INVX1_1/gnd DFFSR_53/S FILL
XINVX1_212 BUFX2_40/Y INVX1_1/gnd INVX1_212/Y DFFSR_97/S INVX1
XFILL_0_INVX1_102 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_1_DFFSR_235 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_7_NAND3X1_35 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_8_OAI22X1_17 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_4_BUFX2_45 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_16_0_0 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_28_DFFSR_162 BUFX2_99/A DFFSR_92/S FILL
XFILL_4_DFFPOSX1_24 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_42_DFFSR_266 INVX1_67/gnd DFFSR_201/S FILL
XFILL_6_NAND3X1_38 BUFX2_98/A DFFSR_32/S FILL
XFILL_4_INVX1_209 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_7_OAI22X1_20 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_18_DFFSR_165 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_32_DFFSR_269 INVX1_67/gnd DFFSR_201/S FILL
XFILL_3_NAND3X1_9 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_6_OAI22X1_23 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_5_NAND3X1_41 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_14_2_1 INVX1_39/gnd DFFSR_54/S FILL
XNAND3X1_38 DFFSR_69/Q BUFX2_16/Y NOR2X1_2/Y BUFX2_98/A NAND3X1_38/Y DFFSR_32/S NAND3X1
XFILL_22_DFFSR_272 INVX1_3/gnd DFFSR_23/S FILL
XFILL_4_NAND3X1_44 BUFX2_99/A DFFSR_7/S FILL
XFILL_9_NAND3X1_139 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_5_OAI22X1_26 INVX1_39/gnd DFFSR_54/S FILL
XFILL_41_DFFSR_67 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_3_NOR2X1_44 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_13_DFFPOSX1_43 OR2X2_2/gnd DFFSR_216/S FILL
XOAI22X1_23 INVX1_54/Y OAI22X1_2/B INVX1_55/Y OAI22X1_2/D DFFSR_4/gnd NOR2X1_27/A
+ DFFSR_4/S OAI22X1
XFILL_12_DFFSR_275 BUFX2_99/A DFFSR_92/S FILL
XFILL_3_NAND3X1_47 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_4_OAI22X1_29 INVX1_3/gnd DFFSR_79/S FILL
XDFFSR_165 DFFSR_165/Q CLKBUF1_10/Y BUFX2_62/Y DFFSR_201/S INVX1_94/A BUFX2_72/gnd
+ DFFSR_201/S DFFSR
XFILL_2_NAND2X1_120 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_12_4_2 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_8_DFFSR_24 BUFX2_98/A DFFSR_6/S FILL
XFILL_2_NAND3X1_50 BUFX2_98/A DFFSR_6/S FILL
XFILL_3_OAI22X1_32 INVX1_39/gnd DFFSR_54/S FILL
XFILL_25_DFFSR_17 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_14_DFFSR_57 BUFX2_79/A DFFSR_6/S FILL
XFILL_4_DFFSR_162 BUFX2_99/A DFFSR_92/S FILL
XFILL_1_BUFX2_92 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_1_NAND3X1_53 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_2_OAI22X1_35 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_45_DFFSR_193 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_8_DFFSR_269 INVX1_67/gnd DFFSR_201/S FILL
XFILL_0_NAND3X1_56 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_1_OAI22X1_38 AND2X2_38/B DFFSR_23/S FILL
XFILL_0_OAI21X1_102 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_35_DFFSR_196 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_23_DFFPOSX1_32 INVX1_67/gnd DFFSR_201/S FILL
XFILL_0_OAI22X1_41 INVX1_39/gnd DFFSR_54/S FILL
XFILL_25_DFFSR_199 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_49_DFFSR_74 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_7_5 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_15_DFFSR_202 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_7_NAND3X1_235 DFFSR_4/gnd DFFSR_4/S FILL
XINVX1_58 INVX1_58/A NOR3X1_6/gnd INVX1_58/Y DFFSR_79/S INVX1
XFILL_33_DFFSR_24 BUFX2_98/A DFFSR_6/S FILL
XFILL_5_DFFSR_71 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_22_DFFSR_64 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_0_NOR2X1_81 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_48_DFFSR_120 INVX1_3/gnd DFFSR_23/S FILL
XFILL_38_DFFSR_123 XOR2X1_4/gnd DFFSR_97/S FILL
XINVX1_176 XNOR2X1_2/Y DFFSR_8/gnd INVX1_176/Y DFFSR_60/S INVX1
XFILL_8_NAND3X1_169 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_1_DFFSR_199 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_28_DFFSR_126 BUFX2_99/A DFFSR_7/S FILL
XFILL_9_XOR2X1_1 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_1_NAND2X1_150 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_42_DFFSR_230 INVX1_67/gnd DFFSR_201/S FILL
XFILL_7_AND2X2_40 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_4_DFFSR_1 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_18_DFFSR_129 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_32_DFFSR_233 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_8_AOI21X1_8 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_22_DFFSR_236 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_9_NAND3X1_103 AND2X2_38/B DFFSR_23/S FILL
XFILL_2_INVX1_65 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_41_DFFSR_31 BUFX2_79/A DFFSR_6/S FILL
XFILL_30_DFFSR_71 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_12_DFFSR_239 INVX1_39/gnd DFFSR_54/S FILL
XFILL_3_NAND3X1_11 OR2X2_4/gnd DFFSR_32/S FILL
XDFFSR_129 DFFSR_153/D CLKBUF1_11/Y BUFX2_67/Y DFFSR_151/S BUFX2_82/A XOR2X1_1/gnd
+ DFFSR_151/S DFFSR
XFILL_2_NAND3X1_14 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_46_1 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_14_DFFSR_21 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_4_DFFSR_126 BUFX2_99/A DFFSR_7/S FILL
XFILL_1_BUFX2_56 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_1_NAND3X1_17 BUFX2_99/A DFFSR_7/S FILL
XFILL_2_OR2X2_1 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_2_0_2 INVX1_67/gnd DFFSR_201/S FILL
XFILL_45_DFFSR_157 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_11_AOI22X1_4 BUFX2_99/A DFFSR_92/S FILL
XFILL_8_DFFSR_233 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_0_NAND3X1_20 BUFX2_99/A DFFSR_7/S FILL
XFILL_5_NOR3X1_2 INVX1_1/gnd DFFSR_53/S FILL
XFILL_35_DFFSR_160 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_49_DFFSR_264 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_28_DFFSR_5 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_25_DFFSR_163 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_38_DFFSR_78 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_49_DFFSR_38 BUFX2_98/A DFFSR_6/S FILL
XFILL_1_INVX1_210 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_39_DFFSR_267 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_7_NAND3X1_199 INVX1_1/gnd DFFSR_97/S FILL
XFILL_15_DFFSR_166 AND2X2_38/B DFFSR_59/S FILL
XFILL_29_DFFSR_270 INVX1_39/gnd DFFSR_54/S FILL
XFILL_3_DFFPOSX1_18 DFFSR_46/gnd DFFSR_62/S FILL
XINVX1_22 INVX1_22/A OR2X2_4/gnd INVX1_22/Y DFFSR_32/S INVX1
XFILL_0_NAND2X1_180 INVX1_1/gnd DFFSR_97/S FILL
XDFFSR_75 DFFSR_75/Q AOI21X1_3/B DFFSR_1/R DFFSR_1/S DFFSR_67/Q DFFSR_34/gnd DFFSR_1/S
+ DFFSR
XFILL_19_DFFSR_273 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_5_DFFSR_35 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_22_DFFSR_28 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_11_DFFSR_68 BUFX2_98/A DFFSR_6/S FILL
XFILL_49_2_0 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_0_NOR2X1_45 DFFSR_34/gnd DFFSR_1/S FILL
XINVX1_140 INVX1_140/A OR2X2_2/gnd AND2X2_30/B DFFSR_175/S INVX1
XFILL_8_NAND3X1_133 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_47_4_1 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_1_DFFSR_163 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_12_DFFPOSX1_37 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_1_NAND2X1_114 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_4_INVX1_137 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_42_DFFSR_194 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_49_DFFSR_1 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_46_DFFSR_85 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_5_DFFSR_270 INVX1_39/gnd DFFSR_54/S FILL
XFILL_32_DFFSR_197 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_45_6_2 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_22_DFFSR_200 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_30_DFFSR_35 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_2_INVX1_29 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_2_DFFSR_82 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_19_DFFSR_75 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_12_DFFSR_203 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_22_DFFPOSX1_26 AND2X2_38/B DFFSR_23/S FILL
XFILL_6_NAND3X1_229 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_1_BUFX2_20 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_45_DFFSR_121 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_2_DFFPOSX1_48 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_14_XNOR2X1_3 INVX1_1/gnd DFFSR_97/S FILL
XFILL_8_DFFSR_197 XOR2X1_4/gnd DFFSR_97/S FILL
XNOR3X1_6 NOR3X1_6/A NOR3X1_6/B NOR3X1_6/C NOR3X1_6/gnd NOR3X1_6/Y DFFSR_79/S NOR3X1
XFILL_35_DFFSR_124 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_49_DFFSR_228 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_13_5_0 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_25_DFFSR_127 BUFX2_99/A DFFSR_92/S FILL
XFILL_1_INVX1_174 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_38_DFFSR_42 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_39_DFFSR_231 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_27_DFFSR_82 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_4_AND2X2_41 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_15_DFFSR_130 BUFX2_79/A DFFSR_6/S FILL
XFILL_7_NAND3X1_163 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_29_DFFSR_234 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_5_AOI21X1_9 XOR2X1_1/gnd DFFSR_151/S FILL
XDFFSR_39 DFFSR_39/Q CLKBUF1_8/Y DFFSR_7/R DFFSR_79/S DFFSR_23/Q INVX1_3/gnd DFFSR_79/S
+ DFFSR
XFILL_19_DFFSR_237 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_0_NAND2X1_144 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_11_DFFSR_32 OR2X2_4/gnd DFFSR_32/S FILL
XINVX1_104 DFFSR_183/Q BUFX2_7/gnd INVX1_104/Y DFFSR_151/S INVX1
XFILL_1_DFFSR_127 BUFX2_99/A DFFSR_92/S FILL
XFILL_42_DFFSR_158 INVX1_3/gnd DFFSR_23/S FILL
XFILL_4_INVX1_101 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_46_DFFSR_49 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_35_DFFSR_89 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_5_DFFSR_234 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_32_DFFSR_161 INVX1_67/gnd DFFSR_175/S FILL
XFILL_46_DFFSR_265 INVX1_67/gnd DFFSR_175/S FILL
XFILL_22_DFFSR_164 OR2X2_2/gnd DFFSR_216/S FILL
XAOI22X1_2 NOR3X1_2/Y DFFSR_98/Q DFFSR_98/D NOR3X1_1/Y DFFSR_4/gnd AOI22X1_2/Y DFFSR_98/S
+ AOI22X1
XFILL_19_DFFSR_39 INVX1_3/gnd DFFSR_79/S FILL
XFILL_36_DFFSR_268 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_2_DFFSR_46 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_7_NAND3X1_8 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_6_BUFX2_74 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_12_DFFSR_167 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_26_DFFSR_271 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_8_OAI21X1_115 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_16_DFFSR_274 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_20_CLKBUF1_29 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_6_NAND3X1_193 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_12_XOR2X1_9 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_23_0_0 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_2_DFFPOSX1_12 AND2X2_38/B DFFSR_23/S FILL
XFILL_19_CLKBUF1_32 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_8_DFFSR_161 INVX1_67/gnd DFFSR_175/S FILL
XFILL_43_DFFSR_96 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_18_CLKBUF1_35 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_49_DFFSR_192 INVX1_1/gnd DFFSR_97/S FILL
XNAND3X1_229 INVX1_177/Y NAND2X1_108/Y OAI21X1_79/Y OR2X2_3/gnd NAND3X1_229/Y DFFSR_4/S
+ NAND3X1
XFILL_4_AND2X2_5 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_21_2_1 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_17_CLKBUF1_38 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_1_INVX1_138 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_39_DFFSR_195 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_16_DFFSR_86 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_27_DFFSR_46 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_7_NAND3X1_127 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_2_DFFSR_271 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_3_1_0 INVX1_67/gnd DFFSR_175/S FILL
XFILL_29_DFFSR_198 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_16_CLKBUF1_41 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_11_DFFPOSX1_31 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_19_DFFSR_201 INVX1_67/gnd DFFSR_201/S FILL
XFILL_0_NAND2X1_108 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_15_CLKBUF1_44 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_19_4_2 DFFSR_1/gnd DFFSR_81/S FILL
XNOR2X1_83 NOR2X1_83/A NOR2X1_83/B OR2X2_6/gnd NOR2X1_83/Y DFFSR_92/S NOR2X1
XFILL_1_3_1 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_14_CLKBUF1_47 BUFX2_98/A DFFSR_32/S FILL
XFILL_4_NOR2X1_80 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_40_DFFSR_8 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_42_DFFSR_122 BUFX2_79/A DFFSR_7/S FILL
XFILL_21_DFFPOSX1_20 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_24_DFFSR_93 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_46_DFFSR_13 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_35_DFFSR_53 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_5_DFFSR_198 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_11_XNOR2X1_4 BUFX2_98/A DFFSR_6/S FILL
XFILL_32_DFFSR_125 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_46_DFFSR_229 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_5_NAND3X1_223 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_22_DFFSR_128 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_2_DFFSR_10 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_1_DFFPOSX1_42 INVX1_39/gnd DFFSR_34/S FILL
XFILL_36_DFFSR_232 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_1_AND2X2_42 INVX1_3/gnd DFFSR_23/S FILL
XFILL_12_DFFSR_131 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_6_BUFX2_38 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_26_DFFSR_235 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_11_3 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_16_DFFSR_238 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_6_NAND3X1_157 INVX1_3/gnd DFFSR_23/S FILL
XFILL_4_INVX1_94 INVX1_67/gnd DFFSR_201/S FILL
XFILL_43_DFFSR_60 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_8_DFFSR_125 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_49_DFFSR_156 OR2X2_2/gnd DFFSR_175/S FILL
XNAND3X1_193 NOR3X1_5/B AOI21X1_26/B AOI21X1_26/A XOR2X1_1/gnd AOI21X1_25/B DFFSR_208/S
+ NAND3X1
XFILL_1_INVX1_102 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_39_DFFSR_159 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_27_DFFSR_10 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_16_DFFSR_50 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_2_DFFSR_235 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_3_BUFX2_85 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_29_DFFSR_162 BUFX2_99/A DFFSR_92/S FILL
XFILL_43_DFFSR_266 INVX1_67/gnd DFFSR_201/S FILL
XFILL_19_DFFSR_165 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_20_DFFPOSX1_50 INVX1_1/gnd DFFSR_53/S FILL
XFILL_33_DFFSR_269 INVX1_67/gnd DFFSR_201/S FILL
XNOR2X1_47 NOR2X1_47/A NOR2X1_47/B AND2X2_38/B NOR2X1_47/Y DFFSR_23/S NOR2X1
XFILL_4_NAND3X1_9 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_14_CLKBUF1_11 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_23_DFFSR_272 INVX1_3/gnd DFFSR_23/S FILL
XFILL_9_0_2 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_4_NOR2X1_44 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_13_CLKBUF1_14 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_13_DFFSR_275 BUFX2_99/A DFFSR_92/S FILL
XFILL_12_CLKBUF1_17 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_7_OAI21X1_109 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_35_DFFSR_17 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_7_DFFSR_64 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_24_DFFSR_57 BUFX2_79/A DFFSR_6/S FILL
XFILL_11_CLKBUF1_20 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_5_DFFSR_162 BUFX2_99/A DFFSR_92/S FILL
XFILL_13_DFFSR_97 INVX1_1/gnd DFFSR_97/S FILL
XFILL_46_DFFSR_193 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_5_NAND3X1_187 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_10_CLKBUF1_23 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_9_DFFSR_269 INVX1_67/gnd DFFSR_201/S FILL
XFILL_36_DFFSR_196 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_9_CLKBUF1_26 INVX1_1/gnd DFFSR_53/S FILL
XFILL_26_DFFSR_199 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_16_DFFSR_202 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_27_DFFSR_2 BUFX2_79/A DFFSR_7/S FILL
XFILL_8_CLKBUF1_29 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_6_NAND3X1_121 INVX1_1/gnd DFFSR_97/S FILL
XFILL_54_4_1 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_7_CLKBUF1_32 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_10_DFFPOSX1_25 BUFX2_79/A DFFSR_6/S FILL
XFILL_43_DFFSR_24 BUFX2_98/A DFFSR_6/S FILL
XFILL_4_INVX1_58 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_32_DFFSR_64 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_6_CLKBUF1_35 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_1_NOR2X1_81 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_49_DFFSR_120 INVX1_3/gnd DFFSR_23/S FILL
XFILL_5_CLKBUF1_38 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_52_6_2 BUFX2_77/gnd DFFSR_98/S FILL
XNAND3X1_157 BUFX2_58/Y AND2X2_33/B NAND2X1_77/A INVX1_3/gnd NAND3X1_158/B DFFSR_23/S
+ NAND3X1
XCLKBUF1_35 BUFX2_2/Y DFFSR_5/gnd DFFSR_82/CLK DFFSR_5/S CLKBUF1
XFILL_39_DFFSR_123 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_16_DFFSR_14 INVX1_1/gnd DFFSR_53/S FILL
XFILL_4_CLKBUF1_41 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_2_DFFSR_199 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_3_BUFX2_49 INVX1_1/gnd DFFSR_97/S FILL
XFILL_29_DFFSR_126 BUFX2_99/A DFFSR_7/S FILL
XFILL_43_DFFSR_230 INVX1_67/gnd DFFSR_201/S FILL
XFILL_3_CLKBUF1_44 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_8_AND2X2_40 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_19_DFFSR_129 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_20_DFFPOSX1_14 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_33_DFFSR_233 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_2_CLKBUF1_47 BUFX2_98/A DFFSR_32/S FILL
XXNOR2X1_2 NOR2X1_71/B XNOR2X1_2/B BUFX2_98/A XNOR2X1_2/Y DFFSR_6/S XNOR2X1
XNOR2X1_11 NOR2X1_11/A NOR2X1_11/B DFFSR_8/gnd NOR2X1_11/Y DFFSR_60/S NOR2X1
XFILL_9_AOI21X1_8 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_23_DFFSR_236 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_4_NAND3X1_217 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_40_DFFSR_71 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_0_DFFPOSX1_36 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_13_DFFSR_239 INVX1_39/gnd DFFSR_54/S FILL
XFILL_20_5_0 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_7_DFFSR_28 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_24_DFFSR_21 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_13_DFFSR_61 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_5_DFFSR_126 BUFX2_99/A DFFSR_7/S FILL
XFILL_0_BUFX2_96 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_46_DFFSR_157 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_5_NAND3X1_151 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_9_DFFSR_233 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_36_DFFSR_160 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_6_NOR2X1_9 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_50_DFFSR_264 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_0_6_0 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_26_DFFSR_163 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_2_INVX1_210 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_40_DFFSR_267 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_48_DFFSR_78 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_16_DFFSR_166 AND2X2_38/B DFFSR_59/S FILL
XFILL_30_DFFSR_270 INVX1_39/gnd DFFSR_54/S FILL
XFILL_20_DFFSR_273 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_19_DFFPOSX1_44 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_32_DFFSR_28 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_21_DFFSR_68 BUFX2_98/A DFFSR_6/S FILL
XFILL_4_DFFSR_75 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_1_NOR2X1_45 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_10_DFFSR_276 BUFX2_72/gnd DFFSR_276/S FILL
XNAND3X1_121 DFFSR_192/D BUFX2_30/Y BUFX2_26/Y INVX1_1/gnd NAND3X1_124/B DFFSR_97/S
+ NAND3X1
XFILL_3_NAND3X1_247 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_2_DFFSR_163 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_3_BUFX2_13 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_8_XOR2X1_5 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_43_DFFSR_194 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_6_OAI21X1_103 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_6_DFFSR_270 INVX1_39/gnd DFFSR_54/S FILL
XFILL_33_DFFSR_197 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_2_CLKBUF1_11 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_23_DFFSR_200 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_1_CLKBUF1_14 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_4_NAND3X1_181 INVX1_39/gnd DFFSR_54/S FILL
XFILL_40_DFFSR_35 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_1_INVX1_69 INVX1_3/gnd DFFSR_23/S FILL
XFILL_30_0_0 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_29_DFFSR_75 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_0_CLKBUF1_17 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_13_DFFSR_203 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_13_DFFSR_25 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_28_2_1 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_0_BUFX2_60 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_46_DFFSR_121 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_5_NAND3X1_115 BUFX2_79/A DFFSR_7/S FILL
XFILL_15_XNOR2X1_3 INVX1_1/gnd DFFSR_97/S FILL
XFILL_9_DFFSR_197 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_36_DFFSR_124 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_4_NOR3X1_6 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_26_4_2 INVX1_3/gnd DFFSR_23/S FILL
XFILL_50_DFFSR_228 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_18_DFFSR_9 BUFX2_79/A DFFSR_6/S FILL
XFILL_26_DFFSR_127 BUFX2_99/A DFFSR_92/S FILL
XFILL_2_INVX1_174 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_40_DFFSR_231 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_8_3_1 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_37_DFFSR_82 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_48_DFFSR_42 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_5_AND2X2_41 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_16_DFFSR_130 BUFX2_79/A DFFSR_6/S FILL
XFILL_30_DFFSR_234 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_6_AOI21X1_9 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_20_DFFSR_237 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_4_DFFSR_39 INVX1_3/gnd DFFSR_79/S FILL
XFILL_6_5_2 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_10_DFFSR_72 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_21_DFFSR_32 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_10_DFFSR_240 INVX1_39/gnd DFFSR_34/S FILL
XFILL_3_NAND3X1_211 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_2_DFFSR_127 BUFX2_99/A DFFSR_92/S FILL
XFILL_14_XOR2X1_2 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_39_DFFSR_5 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_55_3 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_43_DFFSR_158 INVX1_3/gnd DFFSR_23/S FILL
XFILL_45_DFFSR_89 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_6_DFFSR_234 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_33_DFFSR_161 INVX1_67/gnd DFFSR_175/S FILL
XFILL_47_DFFSR_265 INVX1_67/gnd DFFSR_175/S FILL
XFILL_25_DFFPOSX1_2 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_23_DFFSR_164 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_4_NAND3X1_145 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_1_INVX1_33 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_1_DFFSR_86 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_29_DFFSR_39 INVX1_3/gnd DFFSR_79/S FILL
XFILL_37_DFFSR_268 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_24_DFFPOSX1_5 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_18_DFFSR_79 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_13_DFFSR_167 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_8_NAND3X1_8 XOR2X1_4/gnd DFFSR_97/S FILL
XOAI21X1_103 DFFSR_92/S INVX1_201/Y NAND2X1_134/Y OR2X2_6/gnd DFFSR_275/D DFFSR_92/S
+ OAI21X1
XFILL_27_DFFSR_271 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_23_DFFPOSX1_8 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_9_DFFPOSX1_19 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_6_NAND2X1_181 BUFX2_99/A DFFSR_92/S FILL
XFILL_17_DFFSR_274 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_0_BUFX2_24 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_9_DFFSR_161 INVX1_67/gnd DFFSR_175/S FILL
XFILL_10_NOR3X1_3 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_18_DFFPOSX1_38 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_50_DFFSR_192 INVX1_1/gnd DFFSR_97/S FILL
XFILL_2_INVX1_138 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_40_DFFSR_195 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_9_DFFSR_93 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_26_DFFSR_86 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_37_DFFSR_46 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_2_NAND3X1_241 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_3_DFFSR_271 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_30_DFFSR_198 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_20_DFFSR_201 INVX1_67/gnd DFFSR_201/S FILL
XFILL_10_DFFSR_36 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_10_DFFSR_204 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_3_NAND3X1_175 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_5_NOR2X1_80 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_43_DFFSR_122 BUFX2_79/A DFFSR_7/S FILL
XFILL_8_DFFPOSX1_49 BUFX2_99/A DFFSR_92/S FILL
XFILL_45_DFFSR_53 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_6_DFFSR_198 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_34_DFFSR_93 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_12_XNOR2X1_4 BUFX2_98/A DFFSR_6/S FILL
XFILL_33_DFFSR_125 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_47_DFFSR_229 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_4_NAND3X1_109 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_23_DFFSR_128 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_1_DFFSR_50 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_37_DFFSR_232 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_18_DFFSR_43 BUFX2_98/A DFFSR_6/S FILL
XFILL_2_AND2X2_42 INVX1_3/gnd DFFSR_23/S FILL
XFILL_13_DFFSR_131 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_5_BUFX2_78 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_27_DFFSR_235 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_6_NAND2X1_145 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_17_DFFSR_238 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_6_DFFSR_8 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_9_DFFSR_125 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_9_AOI21X1_70 OR2X2_6/gnd DFFSR_92/S FILL
XNAND2X1_181 XOR2X1_15/A XOR2X1_15/B BUFX2_99/A AOI21X1_71/B DFFSR_92/S NAND2X1
XFILL_50_DFFSR_156 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_3_AND2X2_9 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_2_INVX1_102 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_40_DFFSR_159 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_37_DFFSR_10 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_26_DFFSR_50 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_15_DFFSR_90 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_9_DFFSR_57 BUFX2_79/A DFFSR_6/S FILL
XFILL_2_NAND3X1_205 INVX1_1/gnd DFFSR_53/S FILL
XFILL_3_DFFSR_235 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_10_XOR2X1_10 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_30_DFFSR_162 BUFX2_99/A DFFSR_92/S FILL
XFILL_44_DFFSR_266 INVX1_67/gnd DFFSR_201/S FILL
XFILL_20_DFFSR_165 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_34_DFFSR_269 INVX1_67/gnd DFFSR_201/S FILL
XFILL_27_5_0 INVX1_3/gnd DFFSR_79/S FILL
XFILL_5_NAND3X1_9 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_10_DFFSR_168 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_24_DFFSR_272 INVX1_3/gnd DFFSR_23/S FILL
XFILL_3_NAND3X1_139 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_5_NOR2X1_44 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_14_DFFSR_275 BUFX2_99/A DFFSR_92/S FILL
XFILL_8_DFFPOSX1_13 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_13_DFFPOSX1_2 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_7_6_0 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_45_DFFSR_17 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_5_NAND2X1_175 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_34_DFFSR_57 BUFX2_79/A DFFSR_6/S FILL
XFILL_6_DFFSR_162 BUFX2_99/A DFFSR_92/S FILL
XFILL_23_DFFSR_97 INVX1_1/gnd DFFSR_97/S FILL
XFILL_12_DFFPOSX1_5 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_47_DFFSR_193 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_11_DFFPOSX1_8 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_37_DFFSR_196 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_1_DFFSR_14 INVX1_1/gnd DFFSR_53/S FILL
XBUFX2_82 BUFX2_82/A INVX1_1/gnd BUFX2_82/Y DFFSR_97/S BUFX2
XFILL_5_BUFX2_42 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_0_DFFSR_272 INVX1_3/gnd DFFSR_23/S FILL
XFILL_17_DFFPOSX1_32 INVX1_67/gnd DFFSR_201/S FILL
XFILL_27_DFFSR_199 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_6_NAND2X1_109 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_17_DFFSR_202 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_51_DFFSR_8 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_1_NAND3X1_235 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_42_DFFSR_64 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_3_INVX1_98 DFFSR_46/gnd DFFSR_62/S FILL
XNAND2X1_145 DFFSR_208/S DFFPOSX1_34/Q XOR2X1_1/gnd AOI21X1_48/B DFFSR_151/S NAND2X1
XFILL_2_NOR2X1_81 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_50_DFFSR_120 INVX1_3/gnd DFFSR_23/S FILL
XFILL_27_DFFPOSX1_21 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_8_AOI21X1_37 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_40_DFFSR_123 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_9_DFFSR_21 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_26_DFFSR_14 INVX1_1/gnd DFFSR_53/S FILL
XFILL_7_AOI21X1_40 INVX1_39/gnd DFFSR_54/S FILL
XFILL_15_DFFSR_54 INVX1_39/gnd DFFSR_54/S FILL
XFILL_2_NAND3X1_169 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_3_DFFSR_199 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_37_0_0 BUFX2_99/A DFFSR_7/S FILL
XFILL_30_DFFSR_126 BUFX2_99/A DFFSR_7/S FILL
XFILL_2_BUFX2_89 INVX1_1/gnd DFFSR_97/S FILL
XFILL_6_AOI21X1_43 INVX1_3/gnd DFFSR_79/S FILL
XFILL_44_DFFSR_230 INVX1_67/gnd DFFSR_201/S FILL
XFILL_7_DFFPOSX1_43 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_20_DFFSR_129 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_5_AOI21X1_46 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_34_DFFSR_233 OR2X2_2/gnd DFFSR_175/S FILL
XAOI21X1_43 OAI21X1_83/Y INVX1_180/A BUFX2_55/Y INVX1_3/gnd AOI21X1_43/Y DFFSR_79/S
+ AOI21X1
XFILL_35_2_1 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_10_DFFSR_132 INVX1_3/gnd DFFSR_79/S FILL
XFILL_4_AOI21X1_49 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_24_DFFSR_236 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_50_DFFSR_71 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_3_NAND3X1_103 AND2X2_38/B DFFSR_23/S FILL
XFILL_3_AOI21X1_52 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_20_5 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_14_DFFSR_239 INVX1_39/gnd DFFSR_54/S FILL
XFILL_33_4_2 INVX1_1/gnd DFFSR_53/S FILL
XFILL_2_AOI21X1_55 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_34_DFFSR_21 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_6_DFFSR_68 BUFX2_98/A DFFSR_6/S FILL
XFILL_5_NAND2X1_139 INVX1_1/gnd DFFSR_97/S FILL
XFILL_23_DFFSR_61 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_6_DFFSR_126 BUFX2_99/A DFFSR_7/S FILL
XFILL_1_AOI21X1_58 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_47_DFFSR_157 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_0_AOI21X1_61 AND2X2_38/B DFFSR_59/S FILL
XFILL_37_DFFSR_160 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_51_DFFSR_264 DFFSR_4/gnd DFFSR_98/S FILL
XBUFX2_46 INVX1_59/Y BUFX2_98/A DFFSR_2/R DFFSR_6/S BUFX2
XFILL_0_DFFSR_236 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_27_DFFSR_163 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_3_INVX1_210 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_41_DFFSR_267 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_17_DFFSR_166 AND2X2_38/B DFFSR_59/S FILL
XFILL_17_DFFSR_6 BUFX2_79/A DFFSR_6/S FILL
XFILL_31_DFFSR_270 INVX1_39/gnd DFFSR_54/S FILL
XFILL_8_OAI21X1_85 INVX1_39/gnd DFFSR_54/S FILL
XFILL_1_NAND3X1_199 INVX1_1/gnd DFFSR_97/S FILL
XFILL_7_OAI21X1_88 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_21_DFFSR_273 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_42_DFFSR_28 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_31_DFFSR_68 BUFX2_98/A DFFSR_6/S FILL
XFILL_3_INVX1_62 DFFSR_62/gnd DFFSR_62/S FILL
XNAND2X1_109 INVX1_159/A AND2X2_33/B XOR2X1_4/gnd XNOR2X1_3/B DFFSR_91/S NAND2X1
XFILL_2_NOR2X1_45 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_6_OAI21X1_91 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_11_DFFSR_276 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_5_OAI21X1_94 INVX1_67/gnd DFFSR_175/S FILL
XFILL_1_BUFX2_7 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_15_DFFSR_18 NOR3X1_6/gnd DFFSR_91/S FILL
XOAI21X1_91 DFFSR_51/S INVX1_187/Y OAI21X1_91/C BUFX2_8/gnd DFFSR_263/D DFFSR_51/S
+ OAI21X1
XFILL_2_NAND3X1_133 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_3_DFFSR_163 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_4_OAI21X1_97 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_2_BUFX2_53 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_44_DFFSR_194 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_5_AOI21X1_10 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_7_DFFSR_270 INVX1_39/gnd DFFSR_54/S FILL
XFILL_4_NAND2X1_169 INVX1_1/gnd DFFSR_53/S FILL
XFILL_34_DFFSR_197 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_38_DFFSR_2 BUFX2_79/A DFFSR_7/S FILL
XFILL_4_AOI21X1_13 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_24_DFFSR_200 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_50_DFFSR_35 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_39_DFFSR_75 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_3_AOI21X1_16 INVX1_67/gnd DFFSR_175/S FILL
XFILL_14_DFFSR_203 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_16_DFFPOSX1_26 AND2X2_38/B DFFSR_23/S FILL
XFILL_1_DFFPOSX1_2 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_2_AOI21X1_19 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_6_DFFSR_32 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_5_NAND2X1_103 AND2X2_38/B DFFSR_23/S FILL
XFILL_0_DFFPOSX1_5 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_23_DFFSR_25 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_12_DFFSR_65 BUFX2_79/A DFFSR_7/S FILL
XFILL_1_AOI21X1_22 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_0_NAND3X1_229 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_47_DFFSR_121 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_0_AOI21X1_25 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_16_XNOR2X1_3 INVX1_1/gnd DFFSR_97/S FILL
XFILL_37_DFFSR_124 OR2X2_1/gnd DFFSR_59/S FILL
XBUFX2_10 BUFX2_7/A OR2X2_1/gnd OR2X2_1/B DFFSR_59/S BUFX2
XFILL_0_DFFSR_200 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_27_DFFSR_127 BUFX2_99/A DFFSR_92/S FILL
XFILL_26_DFFPOSX1_15 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_3_INVX1_174 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_41_DFFSR_231 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_47_DFFSR_82 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_6_AND2X2_41 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_17_DFFSR_130 BUFX2_79/A DFFSR_6/S FILL
XFILL_31_DFFSR_234 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_8_OAI21X1_49 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_1_NAND3X1_163 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_7_AOI21X1_9 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_6_NAND2X1_70 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_7_OAI21X1_52 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_21_DFFSR_237 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_31_DFFSR_32 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_3_INVX1_26 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_3_DFFSR_79 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_6_DFFPOSX1_37 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_20_DFFSR_72 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_5_NAND2X1_73 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_6_OAI21X1_55 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_11_DFFSR_240 INVX1_39/gnd DFFSR_34/S FILL
XNAND2X1_70 INVX1_155/A AOI21X1_18/A OR2X2_2/gnd XOR2X1_3/A DFFSR_216/S NAND2X1
XFILL_4_NAND2X1_76 INVX1_3/gnd DFFSR_23/S FILL
XFILL_5_OAI21X1_58 INVX1_39/gnd DFFSR_54/S FILL
XOAI21X1_55 AOI21X1_19/Y AOI21X1_18/Y INVX1_156/A DFFSR_62/gnd OAI21X1_55/Y DFFSR_208/S
+ OAI21X1
XFILL_3_DFFSR_127 BUFX2_99/A DFFSR_92/S FILL
XFILL_2_BUFX2_17 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_42_5 BUFX2_98/A DFFSR_32/S FILL
XFILL_4_OAI21X1_61 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_3_NAND2X1_79 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_7_XOR2X1_9 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_44_DFFSR_158 INVX1_3/gnd DFFSR_23/S FILL
XFILL_10_AOI22X1_5 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_3_OAI21X1_64 INVX1_1/gnd DFFSR_53/S FILL
XFILL_2_NAND2X1_82 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_7_DFFSR_234 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_4_NAND2X1_133 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_34_DFFSR_161 INVX1_67/gnd DFFSR_175/S FILL
XFILL_2_OAI21X1_67 INVX1_1/gnd DFFSR_97/S FILL
XFILL_1_NAND2X1_85 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_48_DFFSR_265 INVX1_67/gnd DFFSR_175/S FILL
XFILL_24_DFFSR_164 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_1_OAI21X1_70 INVX1_3/gnd DFFSR_23/S FILL
XFILL_38_DFFSR_268 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_0_NAND2X1_88 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_28_DFFSR_79 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_39_DFFSR_39 INVX1_3/gnd DFFSR_79/S FILL
XFILL_0_INVX1_211 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_0_INVX1_73 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_9_NAND3X1_8 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_14_DFFSR_167 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_0_OAI21X1_73 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_28_DFFSR_271 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_2_OAI21X1_115 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_18_DFFSR_274 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_25_DFFPOSX1_45 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_12_DFFSR_29 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_0_NAND3X1_193 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_9_NAND3X1_248 INVX1_3/gnd DFFSR_79/S FILL
XFILL_5_DFFSR_5 DFFSR_5/gnd DFFSR_5/S FILL
XDFFSR_9 DFFSR_9/Q DFFSR_9/CLK DFFSR_9/R DFFSR_6/S INVX1_1/A BUFX2_79/A DFFSR_6/S
+ DFFSR
XDFFSR_274 BUFX2_72/A CLKBUF1_15/Y DFFSR_274/R DFFSR_276/S DFFSR_274/D BUFX2_72/gnd
+ DFFSR_276/S DFFSR
XFILL_0_DFFSR_164 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_34_5_0 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_3_INVX1_138 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_41_DFFSR_195 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_36_DFFSR_86 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_47_DFFSR_46 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_4_DFFSR_271 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_31_DFFSR_198 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_8_OAI21X1_13 INVX1_39/gnd DFFSR_54/S FILL
XFILL_1_NAND3X1_127 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_7_OAI21X1_16 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_6_NAND2X1_34 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_21_DFFSR_201 INVX1_67/gnd DFFSR_201/S FILL
XFILL_20_DFFSR_36 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_3_DFFSR_43 BUFX2_98/A DFFSR_6/S FILL
XFILL_3_NAND2X1_163 INVX1_67/gnd DFFSR_201/S FILL
XFILL_5_NAND2X1_37 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_6_OAI21X1_19 BUFX2_98/A DFFSR_32/S FILL
XFILL_11_DFFSR_204 BUFX2_7/gnd DFFSR_216/S FILL
XNAND2X1_34 INVX1_62/A NOR3X1_3/A NOR3X1_6/gnd NOR3X1_4/C DFFSR_91/S NAND2X1
XFILL_4_NAND2X1_40 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_3_OR2X2_5 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_6_NOR2X1_80 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_5_OAI21X1_22 DFFSR_34/gnd DFFSR_34/S FILL
XOAI21X1_19 NOR3X1_4/B NOR3X1_4/A AOI21X1_4/Y BUFX2_98/A OAI21X1_19/Y DFFSR_32/S OAI21X1
XFILL_3_NAND2X1_43 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_4_OAI21X1_25 DFFSR_62/gnd DFFSR_62/S FILL
XDFFPOSX1_37 DFFPOSX1_37/Q CLKBUF1_43/Y AOI21X1_47/Y BUFX2_72/gnd DFFSR_201/S DFFPOSX1
XFILL_44_DFFSR_122 BUFX2_79/A DFFSR_7/S FILL
XFILL_13_XOR2X1_6 BUFX2_99/A DFFSR_7/S FILL
XFILL_3_OAI21X1_28 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_29_DFFSR_9 BUFX2_79/A DFFSR_6/S FILL
XFILL_2_NAND2X1_46 INVX1_39/gnd DFFSR_34/S FILL
XFILL_15_DFFPOSX1_20 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_44_DFFSR_93 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_13_XNOR2X1_4 BUFX2_98/A DFFSR_6/S FILL
XFILL_7_DFFSR_198 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_34_DFFSR_125 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_1_NAND2X1_49 INVX1_3/gnd DFFSR_79/S FILL
XFILL_2_OAI21X1_31 AND2X2_38/B DFFSR_23/S FILL
XFILL_48_DFFSR_229 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_24_DFFSR_128 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_5_AND2X2_2 BUFX2_99/A DFFSR_7/S FILL
XFILL_1_OAI21X1_34 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_0_INVX1_37 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_0_NAND2X1_52 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_38_DFFSR_232 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_0_DFFSR_90 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_28_DFFSR_43 BUFX2_98/A DFFSR_6/S FILL
XFILL_0_INVX1_175 BUFX2_99/A DFFSR_7/S FILL
XFILL_17_DFFSR_83 INVX1_3/gnd DFFSR_79/S FILL
XFILL_3_AND2X2_42 INVX1_3/gnd DFFSR_23/S FILL
XFILL_14_DFFSR_131 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_28_DFFSR_235 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_0_OAI21X1_37 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_18_DFFSR_238 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_0_NAND3X1_157 INVX1_3/gnd DFFSR_23/S FILL
XFILL_44_0_0 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_50_DFFSR_5 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_5_DFFPOSX1_31 XOR2X1_4/gnd DFFSR_97/S FILL
XDFFSR_238 DFFSR_238/Q CLKBUF1_25/Y BUFX2_67/Y DFFSR_276/S DFFSR_238/D BUFX2_72/gnd
+ DFFSR_276/S DFFSR
XFILL_0_DFFSR_128 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_6_AOI22X1_12 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_42_2_1 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_3_INVX1_102 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_41_DFFSR_159 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_47_DFFSR_10 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_36_DFFSR_50 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_8_DFFSR_97 INVX1_1/gnd DFFSR_97/S FILL
XFILL_25_DFFSR_90 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_4_DFFSR_235 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_11_XOR2X1_10 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_5_AOI22X1_15 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_31_DFFSR_162 BUFX2_99/A DFFSR_92/S FILL
XAOI22X1_12 NOR3X1_4/Y DFFSR_228/Q DFFSR_220/Q NOR3X1_3/Y XOR2X1_1/gnd AOI22X1_12/Y
+ DFFSR_208/S AOI22X1
XFILL_45_DFFSR_266 INVX1_67/gnd DFFSR_201/S FILL
XFILL_4_AOI22X1_18 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_21_DFFSR_165 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_40_4_2 BUFX2_98/A DFFSR_6/S FILL
XFILL_35_DFFSR_269 INVX1_67/gnd DFFSR_201/S FILL
XFILL_14_DFFPOSX1_50 INVX1_1/gnd DFFSR_53/S FILL
XFILL_3_AOI22X1_21 AND2X2_38/B DFFSR_59/S FILL
XFILL_6_NAND3X1_9 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_3_NAND2X1_127 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_11_DFFSR_168 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_25_DFFSR_272 INVX1_3/gnd DFFSR_23/S FILL
XFILL_2_AOI22X1_24 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_6_NOR2X1_44 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_15_DFFSR_275 BUFX2_99/A DFFSR_92/S FILL
XFILL_11_OAI22X1_45 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_1_AOI22X1_27 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_10_OAI22X1_48 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_2_NAND2X1_10 BUFX2_79/A DFFSR_7/S FILL
XFILL_44_DFFSR_57 BUFX2_79/A DFFSR_6/S FILL
XFILL_33_DFFSR_97 INVX1_1/gnd DFFSR_97/S FILL
XFILL_1_OAI21X1_109 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_24_DFFPOSX1_39 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_7_DFFSR_162 BUFX2_99/A DFFSR_92/S FILL
XFILL_1_NAND2X1_13 BUFX2_99/A DFFSR_92/S FILL
XFILL_48_DFFSR_193 OR2X2_2/gnd DFFSR_175/S FILL
XAND2X2_6 AND2X2_6/A AND2X2_6/B BUFX2_99/A AND2X2_6/Y DFFSR_7/S AND2X2
XFILL_8_NAND3X1_69 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_0_NAND2X1_16 BUFX2_79/A DFFSR_7/S FILL
XFILL_9_OAI22X1_51 INVX1_39/gnd DFFSR_54/S FILL
XFILL_38_DFFSR_196 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_8_NAND3X1_242 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_17_DFFSR_47 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_0_INVX1_139 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_0_DFFSR_54 INVX1_39/gnd DFFSR_54/S FILL
XFILL_2_1 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_4_BUFX2_82 INVX1_1/gnd DFFSR_97/S FILL
XFILL_1_DFFSR_272 INVX1_3/gnd DFFSR_23/S FILL
XFILL_7_NAND3X1_72 INVX1_39/gnd DFFSR_34/S FILL
XFILL_28_DFFSR_199 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_6_NAND3X1_75 BUFX2_79/A DFFSR_7/S FILL
XFILL_18_DFFSR_202 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_5_NAND3X1_78 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_0_NAND3X1_121 INVX1_1/gnd DFFSR_97/S FILL
XNAND3X1_75 BUFX2_91/A AND2X2_16/Y BUFX2_33/Y BUFX2_79/A AND2X2_20/A DFFSR_7/S NAND3X1
XFILL_16_DFFSR_3 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_9_NAND3X1_176 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_4_NAND3X1_81 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_3_NOR2X1_81 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_51_DFFSR_120 INVX1_3/gnd DFFSR_23/S FILL
XFILL_3_NAND3X1_84 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_2_NAND2X1_157 NOR3X1_6/gnd DFFSR_91/S FILL
XDFFSR_202 INVX1_72/A CLKBUF1_12/Y BUFX2_70/Y DFFSR_91/S DFFSR_194/Q NOR3X1_6/gnd
+ DFFSR_91/S DFFSR
XFILL_41_DFFSR_123 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_2_NAND3X1_87 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_8_DFFSR_61 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_36_DFFSR_14 INVX1_1/gnd DFFSR_53/S FILL
XFILL_14_DFFSR_94 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_25_DFFSR_54 INVX1_39/gnd DFFSR_54/S FILL
XFILL_4_DFFSR_199 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_31_DFFSR_126 BUFX2_99/A DFFSR_7/S FILL
XFILL_1_NAND3X1_90 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_45_DFFSR_230 INVX1_67/gnd DFFSR_201/S FILL
XFILL_0_BUFX2_4 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_21_DFFSR_129 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_0_NAND3X1_93 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_35_DFFSR_233 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_14_DFFPOSX1_14 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_11_DFFSR_132 INVX1_3/gnd DFFSR_79/S FILL
XFILL_25_DFFSR_236 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_24_2 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_15_DFFSR_239 INVX1_39/gnd DFFSR_54/S FILL
XFILL_10_OAI22X1_12 DFFSR_28/gnd DFFSR_3/S FILL
XINVX1_95 INVX1_95/A BUFX2_7/gnd INVX1_95/Y DFFSR_216/S INVX1
XFILL_33_DFFSR_61 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_44_DFFSR_21 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_7_DFFSR_126 BUFX2_99/A DFFSR_7/S FILL
XFILL_48_DFFSR_157 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_9_OAI22X1_15 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_8_NAND3X1_33 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_38_DFFSR_160 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_8_NAND3X1_206 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_0_INVX1_103 INVX1_39/gnd DFFSR_54/S FILL
XFILL_0_DFFSR_18 NOR3X1_6/gnd DFFSR_91/S FILL
XINVX1_213 OR2X2_5/Y BUFX2_8/gnd INVX1_213/Y DFFSR_81/S INVX1
XFILL_17_DFFSR_11 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_8_OAI22X1_18 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_7_NAND3X1_36 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_4_BUFX2_46 BUFX2_98/A DFFSR_6/S FILL
XFILL_16_0_1 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_1_DFFSR_236 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_28_DFFSR_163 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_4_DFFPOSX1_25 BUFX2_79/A DFFSR_6/S FILL
XFILL_42_DFFSR_267 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_6_NAND3X1_39 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_7_OAI22X1_21 BUFX2_98/A DFFSR_32/S FILL
XFILL_4_INVX1_210 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_18_DFFSR_166 AND2X2_38/B DFFSR_59/S FILL
XFILL_6_OAI22X1_24 BUFX2_98/A DFFSR_32/S FILL
XFILL_5_NAND3X1_42 BUFX2_79/A DFFSR_6/S FILL
XFILL_32_DFFSR_270 INVX1_39/gnd DFFSR_54/S FILL
XFILL_14_2_2 INVX1_39/gnd DFFSR_54/S FILL
XNAND3X1_39 NAND3X1_37/Y NAND3X1_38/Y AOI22X1_5/Y OR2X2_4/gnd NOR2X1_20/B DFFSR_32/S
+ NAND3X1
XFILL_0_AOI22X1_1 INVX1_1/gnd DFFSR_97/S FILL
XFILL_22_DFFSR_273 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_5_OAI22X1_27 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_4_NAND3X1_45 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_41_DFFSR_68 BUFX2_98/A DFFSR_6/S FILL
XFILL_3_NOR2X1_45 DFFSR_34/gnd DFFSR_1/S FILL
XOAI22X1_24 INVX1_56/Y OAI22X1_6/B INVX1_57/Y OAI22X1_6/D BUFX2_98/A NOR2X1_28/A DFFSR_32/S
+ OAI22X1
XFILL_12_DFFSR_276 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_13_DFFPOSX1_44 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_3_NAND3X1_48 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_4_OAI22X1_30 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_2_NAND2X1_121 OR2X2_4/gnd DFFSR_32/S FILL
XDFFSR_166 DFFSR_174/D CLKBUF1_22/Y BUFX2_61/Y DFFSR_59/S INVX1_101/A AND2X2_38/B
+ DFFSR_59/S DFFSR
XFILL_2_NAND3X1_51 BUFX2_99/A DFFSR_7/S FILL
XFILL_3_OAI22X1_33 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_8_DFFSR_25 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_14_DFFSR_58 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_25_DFFSR_18 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_4_DFFSR_163 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_1_NAND3X1_54 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_1_BUFX2_93 AND2X2_38/B DFFSR_59/S FILL
XFILL_2_OAI22X1_36 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_45_DFFSR_194 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_0_NAND3X1_57 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_1_OAI22X1_39 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_8_DFFSR_270 INVX1_39/gnd DFFSR_54/S FILL
XFILL_35_DFFSR_197 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_0_OAI21X1_103 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_23_DFFPOSX1_33 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_0_OAI22X1_42 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_25_DFFSR_200 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_49_DFFSR_75 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_7_6 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_7_NAND3X1_236 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_15_DFFSR_203 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_41_5_0 BUFX2_98/A DFFSR_32/S FILL
XINVX1_59 BUFX2_35/Y OR2X2_1/gnd INVX1_59/Y DFFSR_59/S INVX1
XFILL_5_DFFSR_72 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_33_DFFSR_25 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_22_DFFSR_65 BUFX2_79/A DFFSR_7/S FILL
XFILL_0_NOR2X1_82 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_48_DFFSR_121 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_38_DFFSR_124 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_8_NAND3X1_170 XOR2X1_1/gnd DFFSR_208/S FILL
XINVX1_177 INVX1_177/A OR2X2_3/gnd INVX1_177/Y DFFSR_60/S INVX1
XFILL_4_BUFX2_10 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_1_DFFSR_200 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_28_DFFSR_127 BUFX2_99/A DFFSR_92/S FILL
XFILL_9_XOR2X1_2 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_1_NAND2X1_151 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_42_DFFSR_231 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_4_INVX1_174 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_4_DFFSR_2 BUFX2_79/A DFFSR_7/S FILL
XFILL_7_AND2X2_41 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_18_DFFSR_130 BUFX2_79/A DFFSR_6/S FILL
XFILL_32_DFFSR_234 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_8_AOI21X1_9 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_22_DFFSR_237 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_2_INVX1_66 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_41_DFFSR_32 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_30_DFFSR_72 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_12_DFFSR_240 INVX1_39/gnd DFFSR_34/S FILL
XFILL_3_NAND3X1_12 OR2X2_4/gnd DFFSR_32/S FILL
XDFFSR_130 DFFSR_154/D CLKBUF1_3/Y BUFX2_63/Y DFFSR_6/S BUFX2_83/A BUFX2_79/A DFFSR_6/S
+ DFFSR
XFILL_2_NAND3X1_15 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_46_2 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_14_DFFSR_22 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_4_DFFSR_127 BUFX2_99/A DFFSR_92/S FILL
XFILL_2_OR2X2_2 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_1_NAND3X1_18 BUFX2_79/A DFFSR_7/S FILL
XFILL_1_BUFX2_57 AND2X2_38/B DFFSR_23/S FILL
XFILL_45_DFFSR_158 INVX1_3/gnd DFFSR_23/S FILL
XFILL_8_DFFSR_234 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_0_NAND3X1_21 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_35_DFFSR_161 INVX1_67/gnd DFFSR_175/S FILL
XFILL_5_NOR3X1_3 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_49_DFFSR_265 INVX1_67/gnd DFFSR_175/S FILL
XFILL_28_DFFSR_6 BUFX2_79/A DFFSR_6/S FILL
XFILL_25_DFFSR_164 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_39_DFFSR_268 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_38_DFFSR_79 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_49_DFFSR_39 INVX1_3/gnd DFFSR_79/S FILL
XFILL_1_INVX1_211 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_51_0_0 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_15_DFFSR_167 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_7_NAND3X1_200 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_29_DFFSR_271 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_3_DFFPOSX1_19 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_19_DFFSR_274 BUFX2_72/gnd DFFSR_276/S FILL
XDFFSR_76 DFFSR_84/D DFFSR_92/CLK DFFSR_2/R DFFSR_7/S DFFSR_76/D BUFX2_79/A DFFSR_7/S
+ DFFSR
XINVX1_23 INVX1_23/A BUFX2_99/A INVX1_23/Y DFFSR_7/S INVX1
XFILL_0_NAND2X1_181 BUFX2_99/A DFFSR_92/S FILL
XFILL_22_DFFSR_29 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_5_DFFSR_36 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_49_2_1 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_11_DFFSR_69 BUFX2_98/A DFFSR_32/S FILL
XFILL_0_NOR2X1_46 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_8_NAND3X1_134 INVX1_39/gnd DFFSR_54/S FILL
XINVX1_141 INVX1_141/A INVX1_67/gnd INVX1_141/Y DFFSR_201/S INVX1
XFILL_47_4_2 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_1_DFFSR_164 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_12_DFFPOSX1_38 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_1_NAND2X1_115 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_49_DFFSR_2 BUFX2_79/A DFFSR_7/S FILL
XFILL_42_DFFSR_195 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_4_INVX1_138 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_46_DFFSR_86 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_5_DFFSR_271 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_32_DFFSR_198 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_22_DFFSR_201 INVX1_67/gnd DFFSR_201/S FILL
XFILL_2_INVX1_30 INVX1_1/gnd DFFSR_53/S FILL
XFILL_2_DFFSR_83 INVX1_3/gnd DFFSR_79/S FILL
XFILL_30_DFFSR_36 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_19_DFFSR_76 BUFX2_79/A DFFSR_7/S FILL
XFILL_12_DFFSR_204 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_22_DFFPOSX1_27 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_6_NAND3X1_230 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_1_BUFX2_21 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_15_3_0 INVX1_39/gnd DFFSR_34/S FILL
XFILL_45_DFFSR_122 BUFX2_79/A DFFSR_7/S FILL
XFILL_2_DFFPOSX1_49 BUFX2_99/A DFFSR_92/S FILL
XFILL_8_DFFSR_198 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_14_XNOR2X1_4 BUFX2_98/A DFFSR_6/S FILL
XFILL_35_DFFSR_125 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_49_DFFSR_229 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_13_5_1 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_25_DFFSR_128 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_39_DFFSR_232 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_38_DFFSR_43 BUFX2_98/A DFFSR_6/S FILL
XFILL_1_INVX1_175 BUFX2_99/A DFFSR_7/S FILL
XFILL_27_DFFSR_83 INVX1_3/gnd DFFSR_79/S FILL
XFILL_4_AND2X2_42 INVX1_3/gnd DFFSR_23/S FILL
XFILL_15_DFFSR_131 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_7_NAND3X1_164 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_29_DFFSR_235 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_19_DFFSR_238 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_0_NAND2X1_145 XOR2X1_1/gnd DFFSR_151/S FILL
XDFFSR_40 DFFSR_40/Q DFFSR_8/CLK DFFSR_2/R DFFSR_3/S DFFSR_24/Q OR2X2_4/gnd DFFSR_3/S
+ DFFSR
XFILL_11_DFFSR_33 BUFX2_98/A DFFSR_32/S FILL
XFILL_0_XNOR2X1_1 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_0_NOR2X1_10 BUFX2_98/A DFFSR_32/S FILL
XINVX1_105 DFFSR_183/D BUFX2_7/gnd INVX1_105/Y DFFSR_151/S INVX1
XFILL_1_DFFSR_128 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_42_DFFSR_159 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_46_DFFSR_50 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_35_DFFSR_90 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_5_DFFSR_235 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_12_XOR2X1_10 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_32_DFFSR_162 BUFX2_99/A DFFSR_92/S FILL
XFILL_46_DFFSR_266 INVX1_67/gnd DFFSR_201/S FILL
XFILL_22_DFFSR_165 BUFX2_72/gnd DFFSR_201/S FILL
XAOI22X1_3 NOR3X1_2/Y DFFSR_99/Q DFFSR_91/Q NOR3X1_1/Y INVX1_1/gnd AOI22X1_3/Y DFFSR_97/S
+ AOI22X1
XFILL_2_DFFSR_47 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_36_DFFSR_269 INVX1_67/gnd DFFSR_201/S FILL
XFILL_19_DFFSR_40 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_7_NAND3X1_9 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_6_BUFX2_75 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_12_DFFSR_168 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_26_DFFSR_272 INVX1_3/gnd DFFSR_23/S FILL
XFILL_8_OAI21X1_116 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_16_DFFSR_275 BUFX2_99/A DFFSR_92/S FILL
XFILL_20_CLKBUF1_30 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_6_NAND3X1_194 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_23_0_1 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_43_DFFSR_97 INVX1_1/gnd DFFSR_97/S FILL
XFILL_19_CLKBUF1_33 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_2_DFFPOSX1_13 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_8_DFFSR_162 BUFX2_99/A DFFSR_92/S FILL
XFILL_49_DFFSR_193 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_18_CLKBUF1_36 NOR3X1_6/gnd DFFSR_79/S FILL
XNAND3X1_230 XOR2X1_7/Y NAND3X1_228/Y NAND3X1_229/Y DFFSR_4/gnd NAND3X1_235/B DFFSR_4/S
+ NAND3X1
XFILL_4_AND2X2_6 BUFX2_99/A DFFSR_7/S FILL
XFILL_39_DFFSR_196 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_17_CLKBUF1_39 INVX1_1/gnd DFFSR_53/S FILL
XFILL_21_2_2 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_27_DFFSR_47 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_1_INVX1_139 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_16_DFFSR_87 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_7_NAND3X1_128 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_2_DFFSR_272 INVX1_3/gnd DFFSR_23/S FILL
XFILL_3_1_1 INVX1_67/gnd DFFSR_175/S FILL
XFILL_16_CLKBUF1_42 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_29_DFFSR_199 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_11_DFFPOSX1_32 INVX1_67/gnd DFFSR_201/S FILL
XFILL_15_CLKBUF1_45 BUFX2_79/A DFFSR_7/S FILL
XFILL_0_NAND2X1_109 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_19_DFFSR_202 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_14_CLKBUF1_48 INVX1_3/gnd DFFSR_79/S FILL
XFILL_1_3_2 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_40_DFFSR_9 BUFX2_79/A DFFSR_6/S FILL
XFILL_4_NOR2X1_81 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_21_DFFPOSX1_21 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_42_DFFSR_123 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_46_DFFSR_14 INVX1_1/gnd DFFSR_53/S FILL
XFILL_24_DFFSR_94 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_35_DFFSR_54 INVX1_39/gnd DFFSR_54/S FILL
XFILL_5_DFFSR_199 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_32_DFFSR_126 BUFX2_99/A DFFSR_7/S FILL
XFILL_46_DFFSR_230 INVX1_67/gnd DFFSR_201/S FILL
XFILL_5_NAND3X1_224 INVX1_39/gnd DFFSR_54/S FILL
XFILL_22_DFFSR_129 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_36_DFFSR_233 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_2_DFFSR_11 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_1_DFFPOSX1_43 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_48_5_0 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_6_BUFX2_39 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_12_DFFSR_132 INVX1_3/gnd DFFSR_79/S FILL
XFILL_26_DFFSR_236 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_11_4 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_16_DFFSR_239 INVX1_39/gnd DFFSR_54/S FILL
XFILL_6_NAND3X1_158 AND2X2_38/B DFFSR_59/S FILL
XFILL_4_INVX1_95 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_43_DFFSR_61 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_8_DFFSR_126 BUFX2_99/A DFFSR_7/S FILL
XFILL_49_DFFSR_157 XOR2X1_1/gnd DFFSR_151/S FILL
XNAND3X1_194 NAND2X1_79/B AOI21X1_25/A AOI21X1_25/B DFFSR_62/gnd NAND2X1_90/B DFFSR_208/S
+ NAND3X1
XFILL_39_DFFSR_160 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_27_DFFSR_11 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_1_INVX1_103 INVX1_39/gnd DFFSR_54/S FILL
XFILL_16_DFFSR_51 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_2_DFFSR_236 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_3_BUFX2_86 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_29_DFFSR_163 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_43_DFFSR_267 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_19_DFFSR_166 AND2X2_38/B DFFSR_59/S FILL
XFILL_33_DFFSR_270 INVX1_39/gnd DFFSR_54/S FILL
XNOR2X1_48 NOR2X1_48/A NOR2X1_48/B INVX1_39/gnd NOR2X1_48/Y DFFSR_34/S NOR2X1
XFILL_14_CLKBUF1_12 AND2X2_38/B DFFSR_23/S FILL
XFILL_1_AOI22X1_1 INVX1_1/gnd DFFSR_97/S FILL
XFILL_23_DFFSR_273 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_13_CLKBUF1_15 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_4_NOR2X1_45 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_13_DFFSR_276 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_12_CLKBUF1_18 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_7_OAI21X1_110 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_7_DFFSR_65 BUFX2_79/A DFFSR_7/S FILL
XFILL_11_CLKBUF1_21 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_24_DFFSR_58 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_13_DFFSR_98 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_35_DFFSR_18 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_5_DFFSR_163 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_5_NAND3X1_188 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_10_CLKBUF1_24 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_46_DFFSR_194 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_9_DFFSR_270 INVX1_39/gnd DFFSR_54/S FILL
XFILL_36_DFFSR_197 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_9_CLKBUF1_27 INVX1_1/gnd DFFSR_97/S FILL
XFILL_26_DFFSR_200 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_8_CLKBUF1_30 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_16_DFFSR_203 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_27_DFFSR_3 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_6_NAND3X1_122 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_54_4_2 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_7_CLKBUF1_33 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_10_DFFPOSX1_26 AND2X2_38/B DFFSR_23/S FILL
XFILL_43_DFFSR_25 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_32_DFFSR_65 BUFX2_79/A DFFSR_7/S FILL
XFILL_4_INVX1_59 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_1_NOR2X1_82 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_6_CLKBUF1_36 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_49_DFFSR_121 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_5_CLKBUF1_39 INVX1_1/gnd DFFSR_53/S FILL
XNAND3X1_158 INVX1_151/A NAND3X1_158/B NAND2X1_78/Y AND2X2_38/B AOI21X1_11/B DFFSR_59/S
+ NAND3X1
XFILL_39_DFFSR_124 OR2X2_1/gnd DFFSR_59/S FILL
XCLKBUF1_36 BUFX2_4/Y NOR3X1_6/gnd DFFSR_83/CLK DFFSR_79/S CLKBUF1
XFILL_16_DFFSR_15 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_4_CLKBUF1_42 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_2_DFFSR_200 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_3_BUFX2_50 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_29_DFFSR_127 BUFX2_99/A DFFSR_92/S FILL
XFILL_43_DFFSR_231 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_3_CLKBUF1_45 BUFX2_79/A DFFSR_7/S FILL
XFILL_20_DFFPOSX1_15 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_8_AND2X2_41 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_19_DFFSR_130 BUFX2_79/A DFFSR_6/S FILL
XFILL_33_DFFSR_234 OR2X2_3/gnd DFFSR_4/S FILL
XXNOR2X1_3 XNOR2X1_3/A XNOR2X1_3/B INVX1_1/gnd XOR2X1_7/A DFFSR_97/S XNOR2X1
XFILL_2_CLKBUF1_48 INVX1_3/gnd DFFSR_79/S FILL
XNOR2X1_12 OAI22X1_8/Y OAI22X1_7/Y XOR2X1_4/gnd NOR2X1_12/Y DFFSR_97/S NOR2X1
XFILL_22_3_0 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_23_DFFSR_237 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_4_NAND3X1_218 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_40_DFFSR_72 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_0_DFFPOSX1_37 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_13_DFFSR_240 INVX1_39/gnd DFFSR_34/S FILL
XFILL_20_5_1 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_7_DFFSR_29 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_24_DFFSR_22 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_13_DFFSR_62 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_5_DFFSR_127 BUFX2_99/A DFFSR_92/S FILL
XFILL_0_BUFX2_97 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_2_4_0 INVX1_67/gnd DFFSR_201/S FILL
XFILL_46_DFFSR_158 INVX1_3/gnd DFFSR_23/S FILL
XFILL_5_NAND3X1_152 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_9_DFFSR_234 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_36_DFFSR_161 INVX1_67/gnd DFFSR_175/S FILL
XFILL_3_INVX1_1 INVX1_1/gnd DFFSR_53/S FILL
XFILL_50_DFFSR_265 INVX1_67/gnd DFFSR_175/S FILL
XFILL_0_6_1 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_26_DFFSR_164 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_48_DFFSR_79 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_40_DFFSR_268 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_2_INVX1_211 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_16_DFFSR_167 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_30_DFFSR_271 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_20_DFFSR_274 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_32_DFFSR_29 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_4_DFFSR_76 BUFX2_79/A DFFSR_7/S FILL
XFILL_4_INVX1_23 BUFX2_99/A DFFSR_7/S FILL
XFILL_21_DFFSR_69 BUFX2_98/A DFFSR_32/S FILL
XFILL_19_DFFPOSX1_45 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_1_NOR2X1_46 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_10_DFFSR_277 BUFX2_72/gnd DFFSR_201/S FILL
XNAND3X1_122 DFFSR_136/Q AND2X2_18/B BUFX2_30/Y XOR2X1_4/gnd AND2X2_26/B DFFSR_97/S
+ NAND3X1
XFILL_3_NAND3X1_248 INVX1_3/gnd DFFSR_79/S FILL
XFILL_2_DFFSR_164 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_3_BUFX2_14 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_8_XOR2X1_6 BUFX2_99/A DFFSR_7/S FILL
XFILL_43_DFFSR_195 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_6_OAI21X1_104 INVX1_67/gnd DFFSR_201/S FILL
XFILL_6_DFFSR_271 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_33_DFFSR_198 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_2_CLKBUF1_12 AND2X2_38/B DFFSR_23/S FILL
XFILL_23_DFFSR_201 INVX1_67/gnd DFFSR_201/S FILL
XFILL_4_NAND3X1_182 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_1_CLKBUF1_15 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_40_DFFSR_36 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_29_DFFSR_76 BUFX2_79/A DFFSR_7/S FILL
XFILL_1_INVX1_70 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_30_0_1 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_13_DFFSR_204 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_0_CLKBUF1_18 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_13_DFFSR_26 BUFX2_79/A DFFSR_6/S FILL
XFILL_28_2_2 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_0_BUFX2_61 AND2X2_38/B DFFSR_59/S FILL
XFILL_46_DFFSR_122 BUFX2_79/A DFFSR_7/S FILL
XFILL_5_NAND3X1_116 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_9_DFFSR_198 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_15_XNOR2X1_4 BUFX2_98/A DFFSR_6/S FILL
XFILL_36_DFFSR_125 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_50_DFFSR_229 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_26_DFFSR_128 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_40_DFFSR_232 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_8_3_2 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_48_DFFSR_43 BUFX2_98/A DFFSR_6/S FILL
XFILL_2_INVX1_175 BUFX2_99/A DFFSR_7/S FILL
XFILL_37_DFFSR_83 INVX1_3/gnd DFFSR_79/S FILL
XFILL_5_AND2X2_42 INVX1_3/gnd DFFSR_23/S FILL
XFILL_16_DFFSR_131 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_30_DFFSR_235 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_20_DFFSR_238 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_4_DFFSR_40 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_21_DFFSR_33 BUFX2_98/A DFFSR_32/S FILL
XFILL_10_DFFSR_73 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_1_XNOR2X1_1 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_1_NOR2X1_10 BUFX2_98/A DFFSR_32/S FILL
XFILL_10_DFFSR_241 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_3_NAND3X1_212 INVX1_39/gnd DFFSR_54/S FILL
XFILL_2_DFFSR_128 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_14_XOR2X1_3 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_43_DFFSR_159 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_55_4 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_39_DFFSR_6 BUFX2_79/A DFFSR_6/S FILL
XFILL_45_DFFSR_90 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_6_DFFSR_235 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_13_XOR2X1_10 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_33_DFFSR_162 BUFX2_99/A DFFSR_92/S FILL
XFILL_47_DFFSR_266 INVX1_67/gnd DFFSR_201/S FILL
XFILL_25_DFFPOSX1_3 INVX1_39/gnd DFFSR_34/S FILL
XFILL_23_DFFSR_165 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_4_NAND3X1_146 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_37_DFFSR_269 INVX1_67/gnd DFFSR_201/S FILL
XFILL_29_DFFSR_40 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_18_DFFSR_80 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_1_DFFSR_87 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_1_INVX1_34 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_8_NAND3X1_9 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_24_DFFPOSX1_6 AND2X2_38/B DFFSR_23/S FILL
XFILL_13_DFFSR_168 OR2X2_6/gnd DFFSR_92/S FILL
XOAI21X1_104 DFFSR_276/S INVX1_202/Y OAI21X1_104/C INVX1_67/gnd DFFSR_276/D DFFSR_201/S
+ OAI21X1
XFILL_27_DFFSR_272 INVX1_3/gnd DFFSR_23/S FILL
XFILL_23_DFFPOSX1_9 INVX1_67/gnd DFFSR_201/S FILL
XFILL_9_DFFPOSX1_20 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_6_NAND2X1_182 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_17_DFFSR_275 BUFX2_99/A DFFSR_92/S FILL
XFILL_0_BUFX2_25 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_9_DFFSR_162 BUFX2_99/A DFFSR_92/S FILL
XFILL_50_DFFSR_193 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_18_DFFPOSX1_39 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_10_NOR3X1_4 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_40_DFFSR_196 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_37_DFFSR_47 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_9_DFFSR_94 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_2_INVX1_139 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_26_DFFSR_87 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_2_NAND3X1_242 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_3_DFFSR_272 INVX1_3/gnd DFFSR_23/S FILL
XFILL_30_DFFSR_199 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_20_DFFSR_202 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_10_DFFSR_37 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_10_DFFSR_205 INVX1_3/gnd DFFSR_79/S FILL
XFILL_5_NOR2X1_81 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_3_NAND3X1_176 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_8_DFFPOSX1_50 INVX1_1/gnd DFFSR_53/S FILL
XFILL_43_DFFSR_123 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_34_DFFSR_94 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_45_DFFSR_54 INVX1_39/gnd DFFSR_54/S FILL
XFILL_6_DFFSR_199 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_33_DFFSR_126 BUFX2_99/A DFFSR_7/S FILL
XFILL_47_DFFSR_230 INVX1_67/gnd DFFSR_201/S FILL
XFILL_23_DFFSR_129 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_4_NAND3X1_110 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_37_DFFSR_233 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_18_DFFSR_44 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_1_DFFSR_51 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_13_DFFSR_132 INVX1_3/gnd DFFSR_79/S FILL
XFILL_5_BUFX2_79 BUFX2_79/A DFFSR_7/S FILL
XFILL_15_1 INVX1_39/gnd DFFSR_54/S FILL
XFILL_27_DFFSR_236 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_6_NAND2X1_146 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_17_DFFSR_239 INVX1_39/gnd DFFSR_54/S FILL
XFILL_6_DFFSR_9 BUFX2_79/A DFFSR_6/S FILL
XFILL_9_DFFSR_126 BUFX2_99/A DFFSR_7/S FILL
XFILL_9_AOI21X1_71 BUFX2_99/A DFFSR_92/S FILL
XNAND2X1_182 INVX1_212/Y NAND2X1_182/B OR2X2_6/gnd NOR2X1_83/B DFFSR_92/S NAND2X1
XFILL_50_DFFSR_157 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_40_DFFSR_160 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_9_DFFSR_58 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_37_DFFSR_11 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_2_INVX1_103 INVX1_39/gnd DFFSR_54/S FILL
XFILL_15_DFFSR_91 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_29_3_0 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_26_DFFSR_51 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_2_NAND3X1_206 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_3_DFFSR_236 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_10_XOR2X1_11 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_30_DFFSR_163 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_44_DFFSR_267 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_20_DFFSR_166 AND2X2_38/B DFFSR_59/S FILL
XFILL_27_5_1 INVX1_3/gnd DFFSR_79/S FILL
XFILL_34_DFFSR_270 INVX1_39/gnd DFFSR_54/S FILL
XFILL_10_DFFSR_169 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_2_AOI22X1_1 INVX1_1/gnd DFFSR_97/S FILL
XFILL_24_DFFSR_273 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_9_4_0 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_3_NAND3X1_140 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_5_NOR2X1_45 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_14_DFFSR_276 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_8_DFFPOSX1_14 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_7_6_1 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_13_DFFPOSX1_3 INVX1_39/gnd DFFSR_34/S FILL
XFILL_34_DFFSR_58 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_5_NAND2X1_176 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_45_DFFSR_18 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_23_DFFSR_98 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_6_DFFSR_163 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_12_DFFPOSX1_6 AND2X2_38/B DFFSR_23/S FILL
XFILL_47_DFFSR_194 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_11_DFFPOSX1_9 INVX1_67/gnd DFFSR_201/S FILL
XFILL_1_DFFSR_15 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_37_DFFSR_197 XOR2X1_4/gnd DFFSR_97/S FILL
XBUFX2_83 BUFX2_83/A BUFX2_79/A BUFX2_83/Y DFFSR_7/S BUFX2
XFILL_5_BUFX2_43 AND2X2_38/B DFFSR_23/S FILL
XFILL_0_DFFSR_273 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_17_DFFPOSX1_33 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_27_DFFSR_200 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_6_NAND2X1_110 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_17_DFFSR_203 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_1_NAND3X1_236 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_42_DFFSR_65 BUFX2_79/A DFFSR_7/S FILL
XFILL_9_AOI21X1_35 INVX1_39/gnd DFFSR_54/S FILL
XFILL_3_INVX1_99 DFFSR_46/gnd DFFSR_62/S FILL
XNAND2X1_146 DFFPOSX1_34/Q INVX1_208/Y BUFX2_7/gnd AOI21X1_49/A DFFSR_151/S NAND2X1
XFILL_2_NOR2X1_82 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_10_CLKBUF1_1 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_50_DFFSR_121 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_8_AOI21X1_38 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_27_DFFPOSX1_22 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_40_DFFSR_124 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_9_DFFSR_22 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_26_DFFSR_15 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_15_DFFSR_55 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_7_AOI21X1_41 INVX1_39/gnd DFFSR_34/S FILL
XFILL_3_DFFSR_200 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_2_NAND3X1_170 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_2_BUFX2_90 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_37_0_1 BUFX2_99/A DFFSR_7/S FILL
XFILL_30_DFFSR_127 BUFX2_99/A DFFSR_92/S FILL
XFILL_6_AOI21X1_44 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_44_DFFSR_231 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_7_DFFPOSX1_44 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_20_DFFSR_130 BUFX2_79/A DFFSR_6/S FILL
XFILL_5_AOI21X1_47 INVX1_67/gnd DFFSR_175/S FILL
XFILL_34_DFFSR_234 OR2X2_3/gnd DFFSR_4/S FILL
XAOI21X1_44 OR2X2_4/Y AOI21X1_44/B INVX1_170/Y DFFSR_28/gnd AOI21X1_44/Y DFFSR_3/S
+ AOI21X1
XFILL_10_DFFSR_133 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_4_AOI21X1_50 INVX1_67/gnd DFFSR_175/S FILL
XFILL_35_2_2 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_24_DFFSR_237 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_50_DFFSR_72 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_3_NAND3X1_104 AND2X2_38/B DFFSR_23/S FILL
XFILL_3_AOI21X1_53 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_20_6 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_14_DFFSR_240 INVX1_39/gnd DFFSR_34/S FILL
XFILL_37_1 BUFX2_99/A DFFSR_92/S FILL
XFILL_2_AOI21X1_56 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_5_NAND2X1_140 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_34_DFFSR_22 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_6_DFFSR_69 BUFX2_98/A DFFSR_32/S FILL
XFILL_23_DFFSR_62 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_6_DFFSR_127 BUFX2_99/A DFFSR_92/S FILL
XFILL_1_AOI21X1_59 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_47_DFFSR_158 INVX1_3/gnd DFFSR_23/S FILL
XFILL_0_AOI21X1_62 INVX1_3/gnd DFFSR_23/S FILL
XFILL_37_DFFSR_161 INVX1_67/gnd DFFSR_175/S FILL
XFILL_51_DFFSR_265 INVX1_67/gnd DFFSR_175/S FILL
XBUFX2_47 INVX1_59/Y OR2X2_3/gnd DFFSR_9/R DFFSR_60/S BUFX2
XFILL_0_DFFSR_237 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_27_DFFSR_164 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_9_OAI21X1_83 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_41_DFFSR_268 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_3_INVX1_211 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_17_DFFSR_167 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_8_OAI21X1_86 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_17_DFFSR_7 BUFX2_79/A DFFSR_7/S FILL
XFILL_1_NAND3X1_200 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_31_DFFSR_271 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_21_DFFSR_274 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_7_OAI21X1_89 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_3_INVX1_63 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_42_DFFSR_29 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_31_DFFSR_69 BUFX2_98/A DFFSR_32/S FILL
XNAND2X1_110 INVX1_145/A NOR3X1_6/gnd NOR3X1_6/gnd XOR2X1_7/B DFFSR_91/S NAND2X1
XFILL_2_NOR2X1_46 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_6_OAI21X1_92 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_11_DFFSR_277 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_5_OAI21X1_95 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_1_BUFX2_8 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_15_DFFSR_19 DFFSR_28/gnd DFFSR_8/S FILL
XOAI21X1_92 DFFSR_260/S INVX1_188/Y OAI21X1_92/C BUFX2_77/gnd DFFSR_264/D DFFSR_98/S
+ OAI21X1
XFILL_3_DFFSR_164 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_2_NAND3X1_134 INVX1_39/gnd DFFSR_54/S FILL
XFILL_2_BUFX2_54 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_4_OAI21X1_98 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_44_DFFSR_195 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_7_DFFSR_271 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_4_NAND2X1_170 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_5_AOI21X1_11 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_34_DFFSR_198 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_38_DFFSR_3 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_4_AOI21X1_14 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_24_DFFSR_201 INVX1_67/gnd DFFSR_201/S FILL
XFILL_50_DFFSR_36 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_39_DFFSR_76 BUFX2_79/A DFFSR_7/S FILL
XFILL_14_DFFSR_204 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_3_AOI21X1_17 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_2_AOI21X1_20 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_16_DFFPOSX1_27 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_1_DFFPOSX1_3 INVX1_39/gnd DFFSR_34/S FILL
XFILL_6_DFFSR_33 BUFX2_98/A DFFSR_32/S FILL
XFILL_23_DFFSR_26 BUFX2_79/A DFFSR_6/S FILL
XFILL_5_NAND2X1_104 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_12_DFFSR_66 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_0_DFFPOSX1_6 AND2X2_38/B DFFSR_23/S FILL
XFILL_1_AOI21X1_23 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_0_NAND3X1_230 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_47_DFFSR_122 BUFX2_79/A DFFSR_7/S FILL
XFILL_0_AOI21X1_26 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_37_DFFSR_125 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_51_DFFSR_229 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_0_DFFSR_201 INVX1_67/gnd DFFSR_201/S FILL
XBUFX2_11 AND2X2_1/Y OR2X2_6/gnd BUFX2_11/Y DFFSR_92/S BUFX2
XFILL_27_DFFSR_128 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_26_DFFPOSX1_16 INVX1_67/gnd DFFSR_175/S FILL
XFILL_3_INVX1_175 BUFX2_99/A DFFSR_7/S FILL
XFILL_41_DFFSR_232 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_47_DFFSR_83 INVX1_3/gnd DFFSR_79/S FILL
XFILL_6_AND2X2_42 INVX1_3/gnd DFFSR_23/S FILL
XFILL_17_DFFSR_131 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_8_OAI21X1_50 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_31_DFFSR_235 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_1_NAND3X1_164 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_21_DFFSR_238 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_6_NAND2X1_71 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_7_OAI21X1_53 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_3_INVX1_27 BUFX2_99/A DFFSR_7/S FILL
XFILL_3_DFFSR_80 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_31_DFFSR_33 BUFX2_98/A DFFSR_32/S FILL
XFILL_20_DFFSR_73 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_2_XNOR2X1_1 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_2_NOR2X1_10 BUFX2_98/A DFFSR_32/S FILL
XFILL_6_DFFPOSX1_38 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_11_DFFSR_241 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_5_NAND2X1_74 AND2X2_38/B DFFSR_59/S FILL
XFILL_6_OAI21X1_56 DFFSR_46/gnd DFFSR_54/S FILL
XNAND2X1_71 AND2X2_35/A AND2X2_35/B DFFSR_34/gnd NAND2X1_71/Y DFFSR_34/S NAND2X1
XFILL_4_NAND2X1_77 AND2X2_38/B DFFSR_23/S FILL
XFILL_5_OAI21X1_59 DFFSR_62/gnd DFFSR_208/S FILL
XOAI21X1_56 OAI21X1_74/A INVX1_163/Y AOI21X1_23/Y DFFSR_46/gnd OAI21X1_56/Y DFFSR_54/S
+ OAI21X1
XFILL_3_DFFSR_128 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_4_OAI21X1_62 INVX1_3/gnd DFFSR_79/S FILL
XFILL_3_NAND2X1_80 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_2_BUFX2_18 BUFX2_98/A DFFSR_32/S FILL
XFILL_44_DFFSR_159 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_10_AOI22X1_6 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_3_OAI21X1_65 INVX1_1/gnd DFFSR_53/S FILL
XFILL_2_NAND2X1_83 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_7_DFFSR_235 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_14_XOR2X1_10 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_4_NAND2X1_134 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_34_DFFSR_162 BUFX2_99/A DFFSR_92/S FILL
XFILL_2_OAI21X1_68 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_1_NAND2X1_86 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_48_DFFSR_266 INVX1_67/gnd DFFSR_201/S FILL
XFILL_24_DFFSR_165 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_1_OAI21X1_71 INVX1_3/gnd DFFSR_79/S FILL
XFILL_0_NAND2X1_89 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_38_DFFSR_269 INVX1_67/gnd DFFSR_201/S FILL
XFILL_39_DFFSR_40 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_0_INVX1_74 BUFX2_99/A DFFSR_92/S FILL
XFILL_0_INVX1_212 INVX1_1/gnd DFFSR_97/S FILL
XFILL_28_DFFSR_80 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_14_DFFSR_168 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_28_DFFSR_272 INVX1_3/gnd DFFSR_23/S FILL
XFILL_0_OAI21X1_74 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_2_OAI21X1_116 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_18_DFFSR_275 BUFX2_99/A DFFSR_92/S FILL
XFILL_25_DFFPOSX1_46 INVX1_39/gnd DFFSR_34/S FILL
XFILL_12_DFFSR_30 BUFX2_98/A DFFSR_32/S FILL
XFILL_36_3_0 BUFX2_99/A DFFSR_92/S FILL
XFILL_0_NAND3X1_194 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_5_DFFSR_6 BUFX2_79/A DFFSR_6/S FILL
XFILL_0_DFFSR_165 BUFX2_72/gnd DFFSR_201/S FILL
XDFFSR_275 BUFX2_73/A DFFSR_2/CLK DFFSR_274/R DFFSR_92/S DFFSR_275/D BUFX2_99/A DFFSR_92/S
+ DFFSR
XFILL_34_5_1 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_41_DFFSR_196 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_3_INVX1_139 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_36_DFFSR_87 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_47_DFFSR_47 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_4_DFFSR_272 INVX1_3/gnd DFFSR_23/S FILL
XFILL_8_OAI21X1_14 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_1_NAND3X1_128 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_31_DFFSR_199 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_6_NAND2X1_35 INVX1_67/gnd DFFSR_201/S FILL
XFILL_21_DFFSR_202 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_7_OAI21X1_17 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_20_DFFSR_37 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_3_DFFSR_44 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_3_NAND2X1_164 INVX1_67/gnd DFFSR_175/S FILL
XFILL_11_DFFSR_205 INVX1_3/gnd DFFSR_79/S FILL
XFILL_6_OAI21X1_20 AND2X2_38/B DFFSR_23/S FILL
XFILL_5_NAND2X1_38 BUFX2_8/gnd DFFSR_81/S FILL
XNAND2X1_35 DFFSR_241/D NOR2X1_34/Y INVX1_67/gnd OAI21X1_9/C DFFSR_201/S NAND2X1
XFILL_3_OR2X2_6 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_5_OAI21X1_23 INVX1_67/gnd DFFSR_201/S FILL
XFILL_4_NAND2X1_41 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_6_NOR2X1_81 XOR2X1_4/gnd DFFSR_97/S FILL
XOAI21X1_20 NOR3X1_4/B NOR3X1_4/A NOR3X1_3/A AND2X2_38/B OAI21X1_20/Y DFFSR_23/S OAI21X1
XFILL_4_OAI21X1_26 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_3_NAND2X1_44 INVX1_39/gnd DFFSR_34/S FILL
XDFFPOSX1_38 BUFX2_58/A CLKBUF1_48/Y NOR2X1_75/Y OR2X2_1/gnd DFFSR_51/S DFFPOSX1
XFILL_44_DFFSR_123 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_13_XOR2X1_7 BUFX2_98/A DFFSR_6/S FILL
XFILL_3_OAI21X1_29 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_15_DFFPOSX1_21 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_44_DFFSR_94 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_2_NAND2X1_47 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_7_DFFSR_199 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_34_DFFSR_126 BUFX2_99/A DFFSR_7/S FILL
XFILL_2_OAI21X1_32 AND2X2_38/B DFFSR_59/S FILL
XFILL_1_NAND2X1_50 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_48_DFFSR_230 INVX1_67/gnd DFFSR_201/S FILL
XFILL_24_DFFSR_129 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_1_OAI21X1_35 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_5_AND2X2_3 INVX1_1/gnd DFFSR_53/S FILL
XFILL_0_NAND2X1_53 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_38_DFFSR_233 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_0_INVX1_176 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_28_DFFSR_44 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_0_DFFSR_91 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_0_INVX1_38 AND2X2_38/B DFFSR_23/S FILL
XFILL_17_DFFSR_84 BUFX2_99/A DFFSR_7/S FILL
XFILL_14_DFFSR_132 INVX1_3/gnd DFFSR_79/S FILL
XFILL_0_OAI21X1_38 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_28_DFFSR_236 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_25_DFFPOSX1_10 INVX1_67/gnd DFFSR_201/S FILL
XFILL_18_DFFSR_239 INVX1_39/gnd DFFSR_54/S FILL
XFILL_0_NAND3X1_158 AND2X2_38/B DFFSR_59/S FILL
XFILL_44_0_1 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_50_DFFSR_6 BUFX2_79/A DFFSR_6/S FILL
XFILL_7_AOI22X1_10 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_5_DFFPOSX1_32 INVX1_67/gnd DFFSR_201/S FILL
XFILL_0_DFFSR_129 XOR2X1_1/gnd DFFSR_151/S FILL
XDFFSR_239 DFFSR_239/Q CLKBUF1_6/Y BUFX2_64/Y DFFSR_54/S DFFSR_231/Q INVX1_39/gnd
+ DFFSR_54/S DFFSR
XFILL_6_AOI22X1_13 AND2X2_38/B DFFSR_23/S FILL
XFILL_42_2_2 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_41_DFFSR_160 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_3_INVX1_103 INVX1_39/gnd DFFSR_54/S FILL
XFILL_8_DFFSR_98 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_25_DFFSR_91 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_36_DFFSR_51 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_47_DFFSR_11 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_5_AOI22X1_16 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_4_DFFSR_236 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_11_XOR2X1_11 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_31_DFFSR_163 DFFSR_1/gnd DFFSR_1/S FILL
XAOI22X1_13 NOR3X1_4/Y DFFSR_237/D DFFSR_229/D NOR3X1_3/Y AND2X2_38/B AOI22X1_13/Y
+ DFFSR_23/S AOI22X1
XFILL_4_AOI22X1_19 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_45_DFFSR_267 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_21_DFFSR_166 AND2X2_38/B DFFSR_59/S FILL
XFILL_35_DFFSR_270 INVX1_39/gnd DFFSR_54/S FILL
XFILL_3_AOI22X1_22 INVX1_3/gnd DFFSR_79/S FILL
XFILL_3_NAND2X1_128 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_11_DFFSR_169 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_3_AOI22X1_1 INVX1_1/gnd DFFSR_97/S FILL
XFILL_25_DFFSR_273 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_2_AOI22X1_25 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_6_NOR2X1_45 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_15_DFFSR_276 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_1_AOI22X1_28 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_10_OAI22X1_49 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_44_DFFSR_58 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_2_NAND2X1_11 BUFX2_98/A DFFSR_6/S FILL
XFILL_10_1_0 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_33_DFFSR_98 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_1_OAI21X1_110 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_7_DFFSR_163 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_24_DFFPOSX1_40 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_1_NAND2X1_14 BUFX2_98/A DFFSR_32/S FILL
XFILL_48_DFFSR_194 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_8_NAND3X1_70 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_9_OAI22X1_52 DFFSR_28/gnd DFFSR_3/S FILL
XAND2X2_7 AND2X2_7/A AND2X2_7/B OR2X2_4/gnd AND2X2_7/Y DFFSR_32/S AND2X2
XFILL_0_NAND2X1_17 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_0_INVX1_140 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_8_NAND3X1_243 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_0_DFFSR_55 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_38_DFFSR_197 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_17_DFFSR_48 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_7_NAND3X1_73 INVX1_1/gnd DFFSR_97/S FILL
XFILL_4_BUFX2_83 BUFX2_79/A DFFSR_7/S FILL
XFILL_1_DFFSR_273 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_28_DFFSR_200 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_6_NAND3X1_76 INVX1_1/gnd DFFSR_53/S FILL
XFILL_18_DFFSR_203 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_5_NAND3X1_79 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_0_NAND3X1_122 XOR2X1_4/gnd DFFSR_97/S FILL
XNAND3X1_76 NAND3X1_76/A NAND3X1_73/Y AND2X2_20/Y INVX1_1/gnd NOR2X1_40/A DFFSR_53/S
+ NAND3X1
XFILL_4_NAND3X1_82 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_16_DFFSR_4 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_3_NOR2X1_82 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_11_CLKBUF1_1 DFFSR_8/gnd DFFSR_8/S FILL
XDFFSR_203 INVX1_79/A DFFSR_1/CLK BUFX2_68/Y DFFSR_54/S DFFSR_195/Q DFFSR_46/gnd DFFSR_54/S
+ DFFSR
XFILL_3_NAND3X1_85 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_2_NAND2X1_158 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_41_DFFSR_124 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_2_NAND3X1_88 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_36_DFFSR_15 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_25_DFFSR_55 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_8_DFFSR_62 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_14_DFFSR_95 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_4_DFFSR_200 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_31_DFFSR_127 BUFX2_99/A DFFSR_92/S FILL
XFILL_1_NAND3X1_91 AND2X2_38/B DFFSR_59/S FILL
XFILL_0_BUFX2_5 AND2X2_38/B DFFSR_59/S FILL
XFILL_45_DFFSR_231 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_21_DFFSR_130 BUFX2_79/A DFFSR_6/S FILL
XFILL_0_NAND3X1_94 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_14_DFFPOSX1_15 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_35_DFFSR_234 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_11_DFFSR_133 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_25_DFFSR_237 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_24_3 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_15_DFFSR_240 INVX1_39/gnd DFFSR_34/S FILL
XFILL_11_OAI22X1_10 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_10_OAI22X1_13 INVX1_1/gnd DFFSR_53/S FILL
XINVX1_96 INVX1_96/A BUFX2_77/gnd INVX1_96/Y DFFSR_98/S INVX1
XFILL_44_DFFSR_22 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_7_DFFSR_127 BUFX2_99/A DFFSR_92/S FILL
XFILL_33_DFFSR_62 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_48_DFFSR_158 INVX1_3/gnd DFFSR_23/S FILL
XFILL_8_NAND3X1_34 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_9_OAI22X1_16 AND2X2_38/B DFFSR_59/S FILL
XFILL_38_DFFSR_161 INVX1_67/gnd DFFSR_175/S FILL
XFILL_0_INVX1_104 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_0_DFFSR_19 DFFSR_28/gnd DFFSR_8/S FILL
XINVX1_214 XOR2X1_11/A XOR2X1_4/gnd NOR2X1_80/A DFFSR_97/S INVX1
XFILL_8_NAND3X1_207 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_17_DFFSR_12 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_7_NAND3X1_37 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_4_BUFX2_47 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_8_OAI22X1_19 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_1_DFFSR_237 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_16_0_2 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_28_DFFSR_164 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_4_DFFPOSX1_26 AND2X2_38/B DFFSR_23/S FILL
XFILL_42_DFFSR_268 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_4_INVX1_211 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_7_OAI22X1_22 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_6_NAND3X1_40 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_18_DFFSR_167 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_32_DFFSR_271 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_5_NAND3X1_43 BUFX2_99/A DFFSR_7/S FILL
XFILL_6_OAI22X1_25 INVX1_39/gnd DFFSR_54/S FILL
XFILL_22_DFFSR_274 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_0_AOI22X1_2 DFFSR_4/gnd DFFSR_98/S FILL
XNAND3X1_40 NOR2X1_18/Y NOR2X1_19/Y NOR2X1_20/Y OR2X2_4/gnd XOR2X1_13/A DFFSR_3/S
+ NAND3X1
XFILL_4_NAND3X1_46 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_5_OAI22X1_28 INVX1_3/gnd DFFSR_23/S FILL
XFILL_41_DFFSR_69 BUFX2_98/A DFFSR_32/S FILL
XFILL_3_NOR2X1_46 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_13_DFFPOSX1_45 OR2X2_1/gnd DFFSR_59/S FILL
XOAI22X1_25 INVX1_60/Y OAI22X1_43/B INVX1_61/Y OAI22X1_43/D INVX1_39/gnd NOR2X1_32/B
+ DFFSR_54/S OAI22X1
XFILL_12_DFFSR_277 BUFX2_72/gnd DFFSR_201/S FILL
XDFFSR_167 DFFSR_175/D CLKBUF1_10/Y BUFX2_64/Y DFFSR_216/S DFFSR_167/D OR2X2_2/gnd
+ DFFSR_216/S DFFSR
XFILL_3_NAND3X1_49 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_4_OAI22X1_31 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_2_NAND2X1_122 INVX1_67/gnd DFFSR_175/S FILL
XFILL_2_NAND3X1_52 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_3_OAI22X1_34 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_25_DFFSR_19 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_8_DFFSR_26 BUFX2_79/A DFFSR_6/S FILL
XFILL_14_DFFSR_59 AND2X2_38/B DFFSR_59/S FILL
XFILL_4_DFFSR_164 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_1_NAND3X1_55 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_2_OAI22X1_37 INVX1_3/gnd DFFSR_23/S FILL
XFILL_1_BUFX2_94 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_45_DFFSR_195 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_0_NAND3X1_58 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_8_DFFSR_271 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_1_OAI22X1_40 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_0_OAI21X1_104 INVX1_67/gnd DFFSR_201/S FILL
XFILL_35_DFFSR_198 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_23_DFFPOSX1_34 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_0_OAI22X1_43 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_25_DFFSR_201 INVX1_67/gnd DFFSR_201/S FILL
XFILL_43_3_0 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_49_DFFSR_76 BUFX2_79/A DFFSR_7/S FILL
XFILL_7_7 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_15_DFFSR_204 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_7_NAND3X1_237 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_41_5_1 BUFX2_98/A DFFSR_32/S FILL
XINVX1_60 INVX1_60/A INVX1_39/gnd INVX1_60/Y DFFSR_34/S INVX1
XFILL_5_DFFSR_73 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_22_DFFSR_66 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_33_DFFSR_26 BUFX2_79/A DFFSR_6/S FILL
XFILL_0_NOR2X1_83 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_48_DFFSR_122 BUFX2_79/A DFFSR_7/S FILL
XINVX1_178 XOR2X1_7/Y DFFSR_4/gnd INVX1_178/Y DFFSR_98/S INVX1
XFILL_38_DFFSR_125 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_8_NAND3X1_171 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_1_DFFSR_201 INVX1_67/gnd DFFSR_201/S FILL
XFILL_4_BUFX2_11 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_9_XOR2X1_3 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_28_DFFSR_128 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_1_NAND2X1_152 INVX1_1/gnd DFFSR_97/S FILL
XFILL_4_INVX1_175 BUFX2_99/A DFFSR_7/S FILL
XFILL_42_DFFSR_232 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_4_DFFSR_3 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_7_AND2X2_42 INVX1_3/gnd DFFSR_23/S FILL
XFILL_18_DFFSR_131 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_32_DFFSR_235 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_22_DFFSR_238 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_4_NAND3X1_10 BUFX2_79/A DFFSR_6/S FILL
XFILL_2_INVX1_67 INVX1_67/gnd DFFSR_201/S FILL
XFILL_41_DFFSR_33 BUFX2_98/A DFFSR_32/S FILL
XFILL_30_DFFSR_73 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_3_XNOR2X1_1 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_3_NOR2X1_10 BUFX2_98/A DFFSR_32/S FILL
XFILL_12_DFFSR_241 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_3_NAND3X1_13 DFFSR_4/gnd DFFSR_4/S FILL
XDFFSR_131 DFFSR_155/D CLKBUF1_27/Y BUFX2_61/Y DFFSR_79/S BUFX2_84/A NOR3X1_6/gnd
+ DFFSR_79/S DFFSR
XFILL_2_NAND3X1_16 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_14_DFFSR_23 AND2X2_38/B DFFSR_23/S FILL
XFILL_46_3 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_4_DFFSR_128 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_2_OR2X2_3 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_1_NAND3X1_19 BUFX2_99/A DFFSR_92/S FILL
XFILL_1_BUFX2_58 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_45_DFFSR_159 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_11_AOI22X1_6 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_8_DFFSR_235 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_0_NAND3X1_22 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_15_XOR2X1_10 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_35_DFFSR_162 BUFX2_99/A DFFSR_92/S FILL
XFILL_5_NOR3X1_4 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_49_DFFSR_266 INVX1_67/gnd DFFSR_201/S FILL
XFILL_28_DFFSR_7 BUFX2_79/A DFFSR_7/S FILL
XFILL_25_DFFSR_165 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_39_DFFSR_269 INVX1_67/gnd DFFSR_201/S FILL
XFILL_49_DFFSR_40 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_1_INVX1_212 INVX1_1/gnd DFFSR_97/S FILL
XFILL_38_DFFSR_80 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_51_0_1 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_15_DFFSR_168 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_7_NAND3X1_201 INVX1_1/gnd DFFSR_53/S FILL
XFILL_29_DFFSR_272 INVX1_3/gnd DFFSR_23/S FILL
XFILL_3_DFFPOSX1_20 DFFSR_46/gnd DFFSR_62/S FILL
XINVX1_24 DFFSR_12/D DFFSR_8/gnd INVX1_24/Y DFFSR_60/S INVX1
XFILL_0_NAND2X1_182 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_5_DFFSR_37 DFFSR_8/gnd DFFSR_60/S FILL
XDFFSR_77 DFFSR_77/Q CLKBUF1_7/Y DFFSR_3/R DFFSR_32/S DFFSR_69/Q BUFX2_98/A DFFSR_32/S
+ DFFSR
XFILL_19_DFFSR_275 BUFX2_99/A DFFSR_92/S FILL
XFILL_11_DFFSR_70 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_22_DFFSR_30 BUFX2_98/A DFFSR_32/S FILL
XFILL_49_2_2 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_0_NOR2X1_47 AND2X2_38/B DFFSR_23/S FILL
XFILL_8_NAND3X1_135 BUFX2_8/gnd DFFSR_81/S FILL
XINVX1_142 AOI21X1_7/B DFFSR_62/gnd AOI21X1_9/C DFFSR_62/S INVX1
XFILL_1_DFFSR_165 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_12_DFFPOSX1_39 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_1_NAND2X1_116 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_42_DFFSR_196 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_49_DFFSR_3 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_4_INVX1_139 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_46_DFFSR_87 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_5_DFFSR_272 INVX1_3/gnd DFFSR_23/S FILL
XFILL_32_DFFSR_199 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_22_DFFSR_202 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_30_DFFSR_37 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_2_DFFSR_84 BUFX2_99/A DFFSR_7/S FILL
XFILL_2_INVX1_31 INVX1_1/gnd DFFSR_53/S FILL
XFILL_19_DFFSR_77 BUFX2_98/A DFFSR_32/S FILL
XFILL_17_1_0 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_12_DFFSR_205 INVX1_3/gnd DFFSR_79/S FILL
XFILL_22_DFFPOSX1_28 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_6_NAND3X1_231 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_15_3_1 INVX1_39/gnd DFFSR_34/S FILL
XFILL_1_BUFX2_22 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_4_INVX1_5 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_45_DFFSR_123 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_2_DFFPOSX1_50 INVX1_1/gnd DFFSR_53/S FILL
XFILL_8_DFFSR_199 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_35_DFFSR_126 BUFX2_99/A DFFSR_7/S FILL
XFILL_11_NOR3X1_1 INVX1_3/gnd DFFSR_79/S FILL
XFILL_49_DFFSR_230 INVX1_67/gnd DFFSR_201/S FILL
XFILL_13_5_2 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_25_DFFSR_129 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_39_DFFSR_233 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_1_INVX1_176 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_38_DFFSR_44 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_27_DFFSR_84 BUFX2_99/A DFFSR_7/S FILL
XFILL_15_DFFSR_132 INVX1_3/gnd DFFSR_79/S FILL
XFILL_7_NAND3X1_165 INVX1_39/gnd DFFSR_34/S FILL
XFILL_29_DFFSR_236 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_0_NAND2X1_146 BUFX2_7/gnd DFFSR_151/S FILL
XDFFSR_41 DFFSR_57/D CLKBUF1_7/Y DFFSR_3/R DFFSR_6/S DFFSR_41/D BUFX2_98/A DFFSR_6/S
+ DFFSR
XFILL_19_DFFSR_239 INVX1_39/gnd DFFSR_54/S FILL
XFILL_0_XNOR2X1_2 BUFX2_98/A DFFSR_6/S FILL
XFILL_11_DFFSR_34 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_0_NOR2X1_11 DFFSR_8/gnd DFFSR_60/S FILL
XINVX1_106 INVX1_106/A INVX1_67/gnd INVX1_106/Y DFFSR_201/S INVX1
XFILL_1_DFFSR_129 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_15_DFFSR_1 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_42_DFFSR_160 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_4_INVX1_103 INVX1_39/gnd DFFSR_54/S FILL
XFILL_35_DFFSR_91 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_46_DFFSR_51 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_12_XOR2X1_11 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_5_DFFSR_236 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_32_DFFSR_163 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_46_DFFSR_267 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_22_DFFSR_166 AND2X2_38/B DFFSR_59/S FILL
XAOI22X1_4 NOR3X1_2/Y DFFSR_100/Q DFFSR_92/Q NOR3X1_1/Y BUFX2_99/A AOI22X1_4/Y DFFSR_92/S
+ AOI22X1
XFILL_2_DFFSR_48 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_36_DFFSR_270 INVX1_39/gnd DFFSR_54/S FILL
XFILL_19_DFFSR_41 BUFX2_98/A DFFSR_6/S FILL
XFILL_6_BUFX2_76 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_12_DFFSR_169 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_4_AOI22X1_1 INVX1_1/gnd DFFSR_97/S FILL
XFILL_26_DFFSR_273 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_8_OAI21X1_117 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_16_DFFSR_276 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_20_CLKBUF1_31 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_6_NAND3X1_195 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_23_0_2 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_19_CLKBUF1_34 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_43_DFFSR_98 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_8_DFFSR_163 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_2_DFFPOSX1_14 DFFSR_62/gnd DFFSR_62/S FILL
XAND2X2_10 AND2X2_10/A AND2X2_10/B DFFSR_8/gnd AND2X2_10/Y DFFSR_8/S AND2X2
XFILL_18_CLKBUF1_37 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_49_DFFSR_194 DFFSR_1/gnd DFFSR_81/S FILL
XNAND3X1_231 NAND3X1_235/B NAND3X1_235/C OR2X2_3/Y DFFSR_4/gnd AOI21X1_36/A DFFSR_98/S
+ NAND3X1
XFILL_4_AND2X2_7 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_1_INVX1_140 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_17_CLKBUF1_40 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_39_DFFSR_197 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_27_DFFSR_48 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_16_DFFSR_88 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_7_NAND3X1_129 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_2_DFFSR_273 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_16_CLKBUF1_43 AND2X2_38/B DFFSR_23/S FILL
XFILL_29_DFFSR_200 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_3_1_2 INVX1_67/gnd DFFSR_175/S FILL
XFILL_11_DFFPOSX1_33 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_15_CLKBUF1_46 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_0_NAND2X1_110 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_19_DFFSR_203 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_14_CLKBUF1_49 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_4_NOR2X1_82 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_12_CLKBUF1_1 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_21_DFFPOSX1_22 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_42_DFFSR_124 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_46_DFFSR_15 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_35_DFFSR_55 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_50_3_0 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_24_DFFSR_95 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_5_DFFSR_200 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_32_DFFSR_127 BUFX2_99/A DFFSR_92/S FILL
XFILL_5_NAND3X1_225 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_46_DFFSR_231 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_22_DFFSR_130 BUFX2_79/A DFFSR_6/S FILL
XFILL_1_DFFPOSX1_44 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_2_DFFSR_12 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_36_DFFSR_234 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_48_5_1 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_12_DFFSR_133 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_6_BUFX2_40 INVX1_1/gnd DFFSR_97/S FILL
XFILL_26_DFFSR_237 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_11_5 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_16_DFFSR_240 INVX1_39/gnd DFFSR_34/S FILL
XFILL_6_NAND3X1_159 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_4_INVX1_96 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_8_DFFSR_127 BUFX2_99/A DFFSR_92/S FILL
XFILL_43_DFFSR_62 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_49_DFFSR_158 INVX1_3/gnd DFFSR_23/S FILL
XNAND3X1_195 INVX1_162/A NAND2X1_90/A NAND2X1_90/B DFFSR_46/gnd INVX1_163/A DFFSR_62/S
+ NAND3X1
XFILL_39_DFFSR_161 INVX1_67/gnd DFFSR_175/S FILL
XFILL_1_INVX1_104 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_27_DFFSR_12 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_16_DFFSR_52 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_3_BUFX2_87 INVX1_1/gnd DFFSR_53/S FILL
XFILL_2_DFFSR_237 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_29_DFFSR_164 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_43_DFFSR_268 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_15_CLKBUF1_10 INVX1_67/gnd DFFSR_201/S FILL
XFILL_19_DFFSR_167 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_33_DFFSR_271 BUFX2_8/gnd DFFSR_81/S FILL
XNOR2X1_49 NOR2X1_49/A NOR2X1_49/B AND2X2_38/B NOR2X1_49/Y DFFSR_59/S NOR2X1
XFILL_14_6_0 INVX1_39/gnd DFFSR_54/S FILL
XFILL_14_CLKBUF1_13 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_23_DFFSR_274 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_1_AOI22X1_2 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_51_DFFSR_69 BUFX2_98/A DFFSR_32/S FILL
XFILL_13_CLKBUF1_16 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_4_NOR2X1_46 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_13_DFFSR_277 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_12_CLKBUF1_19 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_7_OAI21X1_111 AND2X2_38/B DFFSR_59/S FILL
XFILL_35_DFFSR_19 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_7_DFFSR_66 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_5_DFFSR_164 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_13_DFFSR_99 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_24_DFFSR_59 AND2X2_38/B DFFSR_59/S FILL
XFILL_11_CLKBUF1_22 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_10_CLKBUF1_25 INVX1_67/gnd DFFSR_201/S FILL
XFILL_5_NAND3X1_189 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_46_DFFSR_195 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_9_DFFSR_271 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_36_DFFSR_198 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_26_DFFSR_201 INVX1_67/gnd DFFSR_201/S FILL
XFILL_9_CLKBUF1_28 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_8_CLKBUF1_31 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_16_DFFSR_204 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_27_DFFSR_4 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_6_NAND3X1_123 BUFX2_99/A DFFSR_7/S FILL
XFILL_7_CLKBUF1_34 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_10_DFFPOSX1_27 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_32_DFFSR_66 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_43_DFFSR_26 BUFX2_79/A DFFSR_6/S FILL
XFILL_4_INVX1_60 INVX1_39/gnd DFFSR_34/S FILL
XFILL_1_NOR2X1_83 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_6_CLKBUF1_37 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_49_DFFSR_122 BUFX2_79/A DFFSR_7/S FILL
XFILL_5_CLKBUF1_40 OR2X2_6/gnd DFFSR_92/S FILL
XNAND3X1_159 AOI21X1_11/C AOI21X1_11/A AOI21X1_11/B BUFX2_8/gnd OAI21X1_46/C DFFSR_51/S
+ NAND3X1
XCLKBUF1_37 BUFX2_1/Y DFFSR_8/gnd CLKBUF1_37/Y DFFSR_60/S CLKBUF1
XFILL_39_DFFSR_125 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_16_DFFSR_16 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_4_CLKBUF1_43 AND2X2_38/B DFFSR_23/S FILL
XFILL_2_DFFSR_201 INVX1_67/gnd DFFSR_201/S FILL
XFILL_3_BUFX2_51 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_29_DFFSR_128 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_24_1_0 AND2X2_38/B DFFSR_59/S FILL
XFILL_3_CLKBUF1_46 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_43_DFFSR_232 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_8_AND2X2_42 INVX1_3/gnd DFFSR_23/S FILL
XFILL_20_DFFPOSX1_16 INVX1_67/gnd DFFSR_175/S FILL
XFILL_19_DFFSR_131 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_33_DFFSR_235 OR2X2_2/gnd DFFSR_216/S FILL
XXNOR2X1_4 XNOR2X1_4/A XNOR2X1_4/B BUFX2_98/A XNOR2X1_4/Y DFFSR_6/S XNOR2X1
XNOR2X1_13 NOR2X1_13/A NOR2X1_13/B BUFX2_99/A NOR2X1_13/Y DFFSR_92/S NOR2X1
XFILL_2_CLKBUF1_49 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_22_3_1 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_23_DFFSR_238 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_4_NAND3X1_219 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_51_DFFSR_33 BUFX2_98/A DFFSR_32/S FILL
XFILL_40_DFFSR_73 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_4_XNOR2X1_1 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_4_NOR2X1_10 BUFX2_98/A DFFSR_32/S FILL
XFILL_13_DFFSR_241 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_0_DFFPOSX1_38 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_4_2_0 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_20_5_2 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_7_DFFSR_30 BUFX2_98/A DFFSR_32/S FILL
XFILL_13_DFFSR_63 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_5_DFFSR_128 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_24_DFFSR_23 AND2X2_38/B DFFSR_23/S FILL
XFILL_0_BUFX2_98 BUFX2_79/A DFFSR_7/S FILL
XFILL_2_4_1 INVX1_67/gnd DFFSR_201/S FILL
XFILL_46_DFFSR_159 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_5_NAND3X1_153 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_9_DFFSR_235 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_36_DFFSR_162 BUFX2_99/A DFFSR_92/S FILL
XFILL_3_INVX1_2 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_50_DFFSR_266 INVX1_67/gnd DFFSR_201/S FILL
XFILL_0_6_2 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_26_DFFSR_165 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_40_DFFSR_269 INVX1_67/gnd DFFSR_201/S FILL
XFILL_48_DFFSR_80 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_2_INVX1_212 INVX1_1/gnd DFFSR_97/S FILL
XFILL_16_DFFSR_168 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_30_DFFSR_272 INVX1_3/gnd DFFSR_23/S FILL
XFILL_20_DFFSR_275 BUFX2_99/A DFFSR_92/S FILL
XFILL_21_DFFSR_70 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_32_DFFSR_30 BUFX2_98/A DFFSR_32/S FILL
XFILL_4_DFFSR_77 BUFX2_98/A DFFSR_32/S FILL
XFILL_1_NOR2X1_47 AND2X2_38/B DFFSR_23/S FILL
XFILL_19_DFFPOSX1_46 INVX1_39/gnd DFFSR_34/S FILL
XFILL_10_DFFSR_278 XOR2X1_1/gnd DFFSR_151/S FILL
XNAND3X1_123 BUFX2_97/A AND2X2_16/Y BUFX2_33/Y BUFX2_99/A AND2X2_26/A DFFSR_7/S NAND3X1
XFILL_3_NAND3X1_249 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_2_DFFSR_165 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_3_BUFX2_15 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_8_XOR2X1_7 BUFX2_98/A DFFSR_6/S FILL
XFILL_3_CLKBUF1_10 INVX1_67/gnd DFFSR_201/S FILL
XFILL_43_DFFSR_196 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_6_OAI21X1_105 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_6_DFFSR_272 INVX1_3/gnd DFFSR_23/S FILL
XFILL_33_DFFSR_199 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_2_CLKBUF1_13 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_23_DFFSR_202 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_1_CLKBUF1_16 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_4_NAND3X1_183 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_40_DFFSR_37 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_1_INVX1_71 BUFX2_79/A DFFSR_6/S FILL
XFILL_29_DFFSR_77 BUFX2_98/A DFFSR_32/S FILL
XFILL_30_0_2 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_13_DFFSR_205 INVX1_3/gnd DFFSR_79/S FILL
XFILL_0_CLKBUF1_19 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_13_DFFSR_27 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_0_BUFX2_62 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_46_DFFSR_123 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_5_NAND3X1_117 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_9_DFFSR_199 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_36_DFFSR_126 BUFX2_99/A DFFSR_7/S FILL
XFILL_50_DFFSR_230 INVX1_67/gnd DFFSR_201/S FILL
XFILL_26_DFFSR_129 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_40_DFFSR_233 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_2_INVX1_176 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_48_DFFSR_44 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_37_DFFSR_84 BUFX2_99/A DFFSR_7/S FILL
XFILL_16_DFFSR_132 INVX1_3/gnd DFFSR_79/S FILL
XFILL_30_DFFSR_236 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_20_DFFSR_239 INVX1_39/gnd DFFSR_54/S FILL
XFILL_19_DFFPOSX1_10 INVX1_67/gnd DFFSR_201/S FILL
XFILL_1_XNOR2X1_2 BUFX2_98/A DFFSR_6/S FILL
XFILL_4_DFFSR_41 BUFX2_98/A DFFSR_6/S FILL
XFILL_21_DFFSR_34 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_1_NOR2X1_11 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_10_DFFSR_74 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_10_DFFSR_242 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_3_NAND3X1_213 INVX1_39/gnd DFFSR_54/S FILL
XFILL_2_DFFSR_129 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_55_5 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_39_DFFSR_7 BUFX2_79/A DFFSR_7/S FILL
XFILL_14_XOR2X1_4 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_43_DFFSR_160 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_45_DFFSR_91 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_13_XOR2X1_11 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_26_DFFPOSX1_1 INVX1_39/gnd DFFSR_34/S FILL
XFILL_6_DFFSR_236 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_33_DFFSR_163 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_47_DFFSR_267 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_25_DFFPOSX1_4 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_23_DFFSR_166 AND2X2_38/B DFFSR_59/S FILL
XFILL_4_NAND3X1_147 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_1_INVX1_35 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_1_DFFSR_88 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_37_DFFSR_270 INVX1_39/gnd DFFSR_54/S FILL
XFILL_24_DFFPOSX1_7 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_29_DFFSR_41 BUFX2_98/A DFFSR_6/S FILL
XFILL_18_DFFSR_81 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_13_DFFSR_169 DFFSR_62/gnd DFFSR_62/S FILL
XOAI21X1_105 DFFSR_201/S INVX1_203/Y NAND2X1_136/Y BUFX2_72/gnd DFFSR_277/D DFFSR_276/S
+ OAI21X1
XFILL_9_DFFPOSX1_21 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_5_AOI22X1_1 INVX1_1/gnd DFFSR_97/S FILL
XFILL_27_DFFSR_273 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_17_DFFSR_276 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_0_BUFX2_26 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_9_DFFSR_163 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_18_DFFPOSX1_40 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_10_NOR3X1_5 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_50_DFFSR_194 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_21_6_0 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_2_INVX1_140 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_40_DFFSR_197 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_37_DFFSR_48 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_26_DFFSR_88 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_9_DFFSR_95 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_2_NAND3X1_243 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_3_DFFSR_273 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_30_DFFSR_200 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_20_DFFSR_203 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_10_DFFSR_38 BUFX2_98/A DFFSR_6/S FILL
XFILL_10_DFFSR_206 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_5_NOR2X1_82 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_3_NAND3X1_177 AND2X2_38/B DFFSR_59/S FILL
XFILL_13_CLKBUF1_1 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_43_DFFSR_124 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_45_DFFSR_55 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_34_DFFSR_95 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_6_DFFSR_200 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_33_DFFSR_127 BUFX2_99/A DFFSR_92/S FILL
XFILL_47_DFFSR_231 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_23_DFFSR_130 BUFX2_79/A DFFSR_6/S FILL
XFILL_4_NAND3X1_111 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_37_DFFSR_234 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_1_DFFSR_52 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_18_DFFSR_45 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_13_DFFSR_133 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_5_BUFX2_80 BUFX2_79/A DFFSR_6/S FILL
XFILL_15_2 INVX1_39/gnd DFFSR_54/S FILL
XFILL_27_DFFSR_237 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_6_NAND2X1_147 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_17_DFFSR_240 INVX1_39/gnd DFFSR_34/S FILL
XFILL_9_DFFSR_127 BUFX2_99/A DFFSR_92/S FILL
XFILL_31_1_0 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_26_DFFSR_1 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_50_DFFSR_158 INVX1_3/gnd DFFSR_23/S FILL
XFILL_40_DFFSR_161 INVX1_67/gnd DFFSR_175/S FILL
XFILL_2_INVX1_104 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_37_DFFSR_12 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_26_DFFSR_52 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_29_3_1 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_9_DFFSR_59 AND2X2_38/B DFFSR_59/S FILL
XFILL_15_DFFSR_92 BUFX2_99/A DFFSR_92/S FILL
XFILL_2_NAND3X1_207 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_10_XOR2X1_12 INVX1_3/gnd DFFSR_23/S FILL
XFILL_3_DFFSR_237 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_30_DFFSR_164 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_44_DFFSR_268 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_20_DFFSR_167 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_27_5_2 INVX1_3/gnd DFFSR_79/S FILL
XFILL_34_DFFSR_271 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_10_DFFSR_170 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_24_DFFSR_274 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_2_AOI22X1_2 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_9_4_1 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_5_NOR2X1_46 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_3_NAND3X1_141 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_14_DFFSR_277 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_14_DFFPOSX1_1 INVX1_39/gnd DFFSR_34/S FILL
XFILL_8_DFFPOSX1_15 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_13_DFFPOSX1_4 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_7_6_2 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_45_DFFSR_19 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_5_NAND2X1_177 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_23_DFFSR_99 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_34_DFFSR_59 AND2X2_38/B DFFSR_59/S FILL
XFILL_6_DFFSR_164 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_12_DFFPOSX1_7 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_47_DFFSR_195 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_37_DFFSR_198 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_1_DFFSR_16 DFFSR_28/gnd DFFSR_3/S FILL
XBUFX2_84 BUFX2_84/A NOR3X1_6/gnd BUFX2_84/Y DFFSR_91/S BUFX2
XFILL_0_DFFSR_274 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_5_BUFX2_44 INVX1_3/gnd DFFSR_79/S FILL
XFILL_27_DFFSR_201 INVX1_67/gnd DFFSR_201/S FILL
XFILL_17_DFFPOSX1_34 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_6_NAND2X1_111 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_17_DFFSR_204 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_1_NAND3X1_237 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_42_DFFSR_66 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_9_AOI21X1_36 BUFX2_77/gnd DFFSR_98/S FILL
XNAND2X1_147 DFFSR_175/S DFFPOSX1_28/Q OR2X2_2/gnd AOI21X1_49/B DFFSR_216/S NAND2X1
XFILL_2_NOR2X1_83 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_10_CLKBUF1_2 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_50_DFFSR_122 BUFX2_79/A DFFSR_7/S FILL
XFILL_8_AOI21X1_39 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_27_DFFPOSX1_23 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_40_DFFSR_125 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_26_DFFSR_16 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_9_DFFSR_23 AND2X2_38/B DFFSR_23/S FILL
XFILL_7_AOI21X1_42 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_15_DFFSR_56 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_2_NAND3X1_171 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_3_DFFSR_201 INVX1_67/gnd DFFSR_201/S FILL
XFILL_2_BUFX2_91 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_37_0_2 BUFX2_99/A DFFSR_7/S FILL
XFILL_30_DFFSR_128 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_6_AOI21X1_45 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_44_DFFSR_232 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_9_AND2X2_42 INVX1_3/gnd DFFSR_23/S FILL
XFILL_20_DFFSR_131 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_7_DFFPOSX1_45 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_34_DFFSR_235 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_5_AOI21X1_48 DFFSR_62/gnd DFFSR_62/S FILL
XAOI21X1_45 AOI21X1_45/A AOI21X1_45/B INVX1_170/A DFFSR_28/gnd AOI21X1_45/Y DFFSR_3/S
+ AOI21X1
XFILL_10_DFFSR_134 INVX1_1/gnd DFFSR_53/S FILL
XFILL_4_AOI21X1_51 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_24_DFFSR_238 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_5_XNOR2X1_1 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_5_NOR2X1_10 BUFX2_98/A DFFSR_32/S FILL
XFILL_50_DFFSR_73 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_3_NAND3X1_105 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_3_AOI21X1_54 AND2X2_38/B DFFSR_59/S FILL
XFILL_14_DFFSR_241 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_37_2 BUFX2_99/A DFFSR_92/S FILL
XFILL_2_AOI21X1_57 INVX1_67/gnd DFFSR_201/S FILL
XFILL_6_DFFSR_70 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_5_NAND2X1_141 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_23_DFFSR_63 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_34_DFFSR_23 AND2X2_38/B DFFSR_23/S FILL
XFILL_1_AOI21X1_60 BUFX2_79/A DFFSR_7/S FILL
XFILL_6_DFFSR_128 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_47_DFFSR_159 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_0_AOI21X1_63 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_37_DFFSR_162 BUFX2_99/A DFFSR_92/S FILL
XBUFX2_48 INVX1_59/Y AND2X2_38/B DFFSR_73/R DFFSR_59/S BUFX2
XFILL_0_DFFSR_238 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_27_DFFSR_165 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_41_DFFSR_269 INVX1_67/gnd DFFSR_201/S FILL
XFILL_9_OAI21X1_84 BUFX2_98/A DFFSR_6/S FILL
XFILL_3_INVX1_212 INVX1_1/gnd DFFSR_97/S FILL
XFILL_17_DFFSR_168 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_17_DFFSR_8 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_8_OAI21X1_87 BUFX2_79/A DFFSR_7/S FILL
XFILL_1_NAND3X1_201 INVX1_1/gnd DFFSR_53/S FILL
XFILL_31_DFFSR_272 INVX1_3/gnd DFFSR_23/S FILL
XFILL_7_OAI21X1_90 BUFX2_98/A DFFSR_32/S FILL
XFILL_21_DFFSR_275 BUFX2_99/A DFFSR_92/S FILL
XFILL_31_DFFSR_70 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_42_DFFSR_30 BUFX2_98/A DFFSR_32/S FILL
XFILL_3_INVX1_64 DFFSR_46/gnd DFFSR_62/S FILL
XNAND2X1_111 AOI21X1_38/B AOI21X1_38/A DFFSR_8/gnd OR2X2_4/A DFFSR_8/S NAND2X1
XFILL_2_NOR2X1_47 AND2X2_38/B DFFSR_23/S FILL
XFILL_6_OAI21X1_93 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_11_DFFSR_278 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_5_OAI21X1_96 AND2X2_38/B DFFSR_59/S FILL
XFILL_1_BUFX2_9 AND2X2_38/B DFFSR_59/S FILL
XOAI21X1_93 BUFX2_54/Y INVX1_190/Y OAI21X1_93/C OR2X2_2/gnd DFFSR_265/D DFFSR_175/S
+ OAI21X1
XFILL_15_DFFSR_20 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_2_NAND3X1_135 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_3_DFFSR_165 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_4_OAI21X1_99 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_2_BUFX2_55 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_44_DFFSR_196 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_7_DFFSR_272 INVX1_3/gnd DFFSR_23/S FILL
XFILL_4_NAND2X1_171 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_5_AOI21X1_12 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_34_DFFSR_199 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_6_NOR3X1_1 INVX1_3/gnd DFFSR_79/S FILL
XFILL_38_DFFSR_4 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_4_AOI21X1_15 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_24_DFFSR_202 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_50_DFFSR_37 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_39_DFFSR_77 BUFX2_98/A DFFSR_32/S FILL
XFILL_3_AOI21X1_18 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_2_DFFPOSX1_1 INVX1_39/gnd DFFSR_34/S FILL
XFILL_14_DFFSR_205 INVX1_3/gnd DFFSR_79/S FILL
XFILL_2_AOI21X1_21 INVX1_39/gnd DFFSR_54/S FILL
XFILL_1_DFFPOSX1_4 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_16_DFFPOSX1_28 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_5_NAND2X1_105 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_6_DFFSR_34 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_23_DFFSR_27 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_0_DFFPOSX1_7 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_28_6_0 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_12_DFFSR_67 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_1_AOI21X1_24 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_0_NAND3X1_231 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_47_DFFSR_123 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_0_AOI21X1_27 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_37_DFFSR_126 BUFX2_99/A DFFSR_7/S FILL
XBUFX2_12 AND2X2_1/Y DFFSR_28/gnd BUFX2_12/Y DFFSR_8/S BUFX2
XFILL_0_DFFSR_202 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_27_DFFSR_129 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_41_DFFSR_233 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_26_DFFPOSX1_17 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_3_INVX1_176 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_47_DFFSR_84 BUFX2_99/A DFFSR_7/S FILL
XFILL_17_DFFSR_132 INVX1_3/gnd DFFSR_79/S FILL
XFILL_8_OAI21X1_51 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_1_NAND3X1_165 INVX1_39/gnd DFFSR_34/S FILL
XFILL_31_DFFSR_236 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_6_NAND2X1_72 AND2X2_38/B DFFSR_59/S FILL
XFILL_7_OAI21X1_54 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_21_DFFSR_239 INVX1_39/gnd DFFSR_54/S FILL
XFILL_3_INVX1_28 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_2_XNOR2X1_2 BUFX2_98/A DFFSR_6/S FILL
XFILL_3_DFFSR_81 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_31_DFFSR_34 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_6_DFFPOSX1_39 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_20_DFFSR_74 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_2_NOR2X1_11 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_5_NAND2X1_75 INVX1_3/gnd DFFSR_79/S FILL
XFILL_11_DFFSR_242 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_6_OAI21X1_57 DFFSR_34/gnd DFFSR_34/S FILL
XNAND2X1_72 AND2X2_35/A INVX1_159/A AND2X2_38/B OAI21X1_36/C DFFSR_59/S NAND2X1
XFILL_4_NAND2X1_78 AND2X2_38/B DFFSR_23/S FILL
XFILL_5_OAI21X1_60 OR2X2_1/gnd DFFSR_51/S FILL
XOAI21X1_57 INVX1_131/Y NAND2X1_90/Y OAI21X1_57/C DFFSR_34/gnd OAI21X1_57/Y DFFSR_34/S
+ OAI21X1
XFILL_3_DFFSR_129 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_4_OAI21X1_63 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_3_NAND2X1_81 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_2_BUFX2_19 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_44_DFFSR_160 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_10_AOI22X1_7 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_3_OAI21X1_66 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_2_NAND2X1_84 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_14_XOR2X1_11 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_7_DFFSR_236 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_34_DFFSR_163 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_4_NAND2X1_135 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_1_NAND2X1_87 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_2_OAI21X1_69 INVX1_3/gnd DFFSR_23/S FILL
XFILL_48_DFFSR_267 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_24_DFFSR_166 AND2X2_38/B DFFSR_59/S FILL
XFILL_1_OAI21X1_72 INVX1_3/gnd DFFSR_23/S FILL
XFILL_38_DFFSR_270 INVX1_39/gnd DFFSR_54/S FILL
XFILL_0_NAND2X1_90 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_39_DFFSR_41 BUFX2_98/A DFFSR_6/S FILL
XFILL_0_INVX1_75 BUFX2_98/A DFFSR_6/S FILL
XFILL_0_INVX1_213 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_28_DFFSR_81 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_38_1_0 BUFX2_79/A DFFSR_7/S FILL
XFILL_14_DFFSR_169 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_0_OAI21X1_75 INVX1_39/gnd DFFSR_54/S FILL
XFILL_6_AOI22X1_1 INVX1_1/gnd DFFSR_97/S FILL
XFILL_28_DFFSR_273 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_2_OAI21X1_117 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_18_DFFSR_276 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_25_DFFPOSX1_47 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_12_DFFSR_31 BUFX2_79/A DFFSR_6/S FILL
XFILL_36_3_1 BUFX2_99/A DFFSR_92/S FILL
XFILL_0_NAND3X1_195 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_5_DFFSR_7 BUFX2_79/A DFFSR_7/S FILL
XFILL_51_DFFSR_194 DFFSR_1/gnd DFFSR_81/S FILL
XDFFSR_276 BUFX2_74/A CLKBUF1_15/Y DFFSR_274/R DFFSR_276/S DFFSR_276/D BUFX2_72/gnd
+ DFFSR_276/S DFFSR
XFILL_0_DFFSR_166 AND2X2_38/B DFFSR_59/S FILL
XFILL_34_5_2 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_41_DFFSR_197 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_9_OAI21X1_12 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_3_INVX1_140 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_47_DFFSR_48 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_36_DFFSR_88 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_4_DFFSR_273 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_8_OAI21X1_15 INVX1_3/gnd DFFSR_79/S FILL
XFILL_31_DFFSR_200 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_1_NAND3X1_129 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_6_NAND2X1_36 INVX1_3/gnd DFFSR_79/S FILL
XFILL_7_OAI21X1_18 INVX1_39/gnd DFFSR_34/S FILL
XFILL_21_DFFSR_203 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_3_DFFSR_45 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_20_DFFSR_38 BUFX2_98/A DFFSR_6/S FILL
XFILL_5_NAND2X1_39 BUFX2_98/A DFFSR_6/S FILL
XFILL_6_OAI21X1_21 AND2X2_38/B DFFSR_59/S FILL
XFILL_11_DFFSR_206 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_3_NAND2X1_165 DFFSR_62/gnd DFFSR_208/S FILL
XNAND2X1_36 AND2X2_16/Y NOR2X1_30/Y INVX1_3/gnd OAI21X1_9/B DFFSR_79/S NAND2X1
XFILL_5_OAI21X1_24 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_4_NAND2X1_42 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_6_NOR2X1_82 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_14_CLKBUF1_1 DFFSR_8/gnd DFFSR_8/S FILL
XOAI21X1_21 BUFX2_9/Y OR2X2_1/A INVX1_129/Y AND2X2_38/B NOR2X1_63/B DFFSR_59/S OAI21X1
XFILL_4_OAI21X1_27 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_3_NAND2X1_45 INVX1_39/gnd DFFSR_34/S FILL
XDFFPOSX1_39 INVX1_135/A CLKBUF1_44/Y AOI21X1_61/Y BUFX2_7/gnd DFFSR_151/S DFFPOSX1
XFILL_13_XOR2X1_8 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_44_DFFSR_124 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_2_NAND2X1_48 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_3_OAI21X1_30 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_15_DFFPOSX1_22 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_44_DFFSR_95 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_7_DFFSR_200 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_34_DFFSR_127 BUFX2_99/A DFFSR_92/S FILL
XFILL_1_NAND2X1_51 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_2_OAI21X1_33 INVX1_3/gnd DFFSR_79/S FILL
XFILL_48_DFFSR_231 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_24_DFFSR_130 BUFX2_79/A DFFSR_6/S FILL
XFILL_5_AND2X2_4 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_38_DFFSR_234 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_0_NAND2X1_54 AND2X2_38/B DFFSR_59/S FILL
XFILL_1_OAI21X1_36 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_17_DFFSR_85 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_28_DFFSR_45 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_0_INVX1_177 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_0_DFFSR_92 BUFX2_99/A DFFSR_92/S FILL
XFILL_0_INVX1_39 INVX1_39/gnd DFFSR_34/S FILL
XFILL_14_DFFSR_133 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_0_OAI21X1_39 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_28_DFFSR_237 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_25_DFFPOSX1_11 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_18_DFFSR_240 INVX1_39/gnd DFFSR_34/S FILL
XFILL_0_NAND3X1_159 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_44_0_2 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_9_NAND3X1_214 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_7_AOI22X1_11 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_50_DFFSR_7 BUFX2_79/A DFFSR_7/S FILL
XFILL_5_DFFPOSX1_33 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_51_DFFSR_158 INVX1_3/gnd DFFSR_23/S FILL
XFILL_0_DFFSR_130 BUFX2_79/A DFFSR_6/S FILL
XDFFSR_240 DFFSR_240/Q CLKBUF1_6/Y BUFX2_66/Y DFFSR_34/S DFFSR_232/Q INVX1_39/gnd
+ DFFSR_34/S DFFSR
XFILL_6_AOI22X1_14 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_41_DFFSR_161 INVX1_67/gnd DFFSR_175/S FILL
XFILL_3_INVX1_104 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_47_DFFSR_12 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_8_DFFSR_99 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_36_DFFSR_52 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_25_DFFSR_92 BUFX2_99/A DFFSR_92/S FILL
XFILL_5_AOI22X1_17 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_11_XOR2X1_12 INVX1_3/gnd DFFSR_23/S FILL
XFILL_4_DFFSR_237 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_31_DFFSR_164 OR2X2_2/gnd DFFSR_216/S FILL
XAOI22X1_14 NOR3X1_4/Y DFFSR_238/D DFFSR_222/Q NOR3X1_3/Y OR2X2_2/gnd AOI22X1_14/Y
+ DFFSR_216/S AOI22X1
XFILL_45_DFFSR_268 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_4_AOI22X1_20 INVX1_39/gnd DFFSR_34/S FILL
XFILL_21_DFFSR_167 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_35_DFFSR_271 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_3_AOI22X1_23 INVX1_39/gnd DFFSR_34/S FILL
XFILL_11_DFFSR_170 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_3_NAND2X1_129 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_25_DFFSR_274 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_3_AOI22X1_2 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_2_AOI22X1_26 INVX1_1/gnd DFFSR_97/S FILL
XFILL_6_NOR2X1_46 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_15_DFFSR_277 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_1_AOI22X1_29 INVX1_1/gnd DFFSR_53/S FILL
XFILL_10_OAI22X1_50 INVX1_3/gnd DFFSR_23/S FILL
XFILL_2_NAND2X1_12 INVX1_3/gnd DFFSR_79/S FILL
XFILL_33_DFFSR_99 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_1_OAI21X1_111 AND2X2_38/B DFFSR_59/S FILL
XFILL_44_DFFSR_59 AND2X2_38/B DFFSR_59/S FILL
XFILL_10_1_1 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_7_DFFSR_164 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_24_DFFPOSX1_41 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_1_NAND2X1_15 BUFX2_99/A DFFSR_92/S FILL
XFILL_48_DFFSR_195 DFFSR_46/gnd DFFSR_62/S FILL
XAND2X2_8 AND2X2_8/A AND2X2_8/B BUFX2_99/A AND2X2_8/Y DFFSR_7/S AND2X2
XFILL_8_NAND3X1_71 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_38_DFFSR_198 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_0_NAND2X1_18 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_0_INVX1_141 INVX1_67/gnd DFFSR_201/S FILL
XFILL_0_DFFSR_56 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_8_NAND3X1_244 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_17_DFFSR_49 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_1_DFFSR_274 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_7_NAND3X1_74 INVX1_1/gnd DFFSR_97/S FILL
XFILL_4_BUFX2_84 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_28_DFFSR_201 INVX1_67/gnd DFFSR_201/S FILL
XFILL_6_NAND3X1_77 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_18_DFFSR_204 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_5_NAND3X1_80 NOR3X1_6/gnd DFFSR_91/S FILL
XNAND3X1_77 DFFSR_194/D BUFX2_31/Y BUFX2_24/Y DFFSR_5/gnd NAND3X1_79/A DFFSR_5/S NAND3X1
XFILL_0_NAND3X1_123 BUFX2_99/A DFFSR_7/S FILL
XFILL_4_NAND3X1_83 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_16_DFFSR_5 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_9_NAND3X1_178 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_3_NOR2X1_83 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_11_CLKBUF1_2 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_3_NAND3X1_86 DFFSR_62/gnd DFFSR_62/S FILL
XDFFSR_204 INVX1_86/A CLKBUF1_15/Y BUFX2_60/Y DFFSR_216/S DFFSR_204/D BUFX2_7/gnd
+ DFFSR_216/S DFFSR
XFILL_2_NAND2X1_159 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_41_DFFSR_125 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_2_NAND3X1_89 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_36_DFFSR_16 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_8_DFFSR_63 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_25_DFFSR_56 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_14_DFFSR_96 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_4_DFFSR_201 INVX1_67/gnd DFFSR_201/S FILL
XFILL_31_DFFSR_128 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_1_NAND3X1_92 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_45_DFFSR_232 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_0_BUFX2_6 BUFX2_79/A DFFSR_6/S FILL
XFILL_21_DFFSR_131 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_0_NAND3X1_95 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_14_DFFPOSX1_16 INVX1_67/gnd DFFSR_175/S FILL
XFILL_35_DFFSR_235 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_35_6_0 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_11_DFFSR_134 INVX1_1/gnd DFFSR_53/S FILL
XFILL_25_DFFSR_238 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_6_XNOR2X1_1 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_6_NOR2X1_10 BUFX2_98/A DFFSR_32/S FILL
XFILL_24_4 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_15_DFFSR_241 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_11_OAI22X1_11 BUFX2_99/A DFFSR_92/S FILL
XFILL_37_DFFSR_1 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_10_OAI22X1_14 OR2X2_4/gnd DFFSR_3/S FILL
XINVX1_97 INVX1_97/A DFFSR_46/gnd INVX1_97/Y DFFSR_62/S INVX1
XFILL_33_DFFSR_63 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_44_DFFSR_23 AND2X2_38/B DFFSR_23/S FILL
XFILL_7_DFFSR_128 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_48_DFFSR_159 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_8_NAND3X1_35 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_9_OAI22X1_17 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_38_DFFSR_162 BUFX2_99/A DFFSR_92/S FILL
XFILL_0_INVX1_105 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_0_DFFSR_20 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_17_DFFSR_13 OR2X2_6/gnd DFFSR_53/S FILL
XINVX1_215 INVX1_215/A NOR3X1_6/gnd NOR2X1_80/B DFFSR_91/S INVX1
XFILL_8_NAND3X1_208 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_1_DFFSR_238 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_8_OAI22X1_20 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_7_NAND3X1_38 BUFX2_98/A DFFSR_32/S FILL
XFILL_4_BUFX2_48 AND2X2_38/B DFFSR_59/S FILL
XFILL_28_DFFSR_165 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_4_DFFPOSX1_27 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_42_DFFSR_269 INVX1_67/gnd DFFSR_201/S FILL
XFILL_7_OAI22X1_23 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_6_NAND3X1_41 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_18_DFFSR_168 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_32_DFFSR_272 INVX1_3/gnd DFFSR_23/S FILL
XXOR2X1_10 XOR2X1_10/A XOR2X1_10/B OR2X2_1/gnd XOR2X1_10/Y DFFSR_59/S XOR2X1
XFILL_5_NAND3X1_44 BUFX2_99/A DFFSR_7/S FILL
XFILL_6_OAI22X1_26 INVX1_39/gnd DFFSR_54/S FILL
XNAND3X1_41 DFFSR_62/D BUFX2_18/Y BUFX2_11/Y OR2X2_6/gnd NAND3X1_41/Y DFFSR_92/S NAND3X1
XFILL_22_DFFSR_275 BUFX2_99/A DFFSR_92/S FILL
XFILL_0_AOI22X1_3 INVX1_1/gnd DFFSR_97/S FILL
XFILL_9_NAND3X1_142 INVX1_67/gnd DFFSR_175/S FILL
XFILL_4_NAND3X1_47 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_5_OAI22X1_29 INVX1_3/gnd DFFSR_79/S FILL
XFILL_41_DFFSR_70 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_3_NOR2X1_47 AND2X2_38/B DFFSR_23/S FILL
XFILL_13_DFFPOSX1_46 INVX1_39/gnd DFFSR_34/S FILL
XOAI22X1_26 INVX1_64/Y OAI22X1_41/B INVX1_65/Y OAI22X1_41/D INVX1_39/gnd NOR2X1_32/A
+ DFFSR_54/S OAI22X1
XFILL_12_DFFSR_278 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_3_NAND3X1_50 BUFX2_98/A DFFSR_6/S FILL
XFILL_4_OAI22X1_32 INVX1_39/gnd DFFSR_54/S FILL
XFILL_2_NAND2X1_123 BUFX2_77/gnd DFFSR_98/S FILL
XDFFSR_168 DFFSR_176/D CLKBUF1_39/Y BUFX2_63/Y DFFSR_92/S INVX1_115/A OR2X2_6/gnd
+ DFFSR_92/S DFFSR
XFILL_2_NAND3X1_53 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_8_DFFSR_27 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_3_OAI22X1_35 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_14_DFFSR_60 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_25_DFFSR_20 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_4_DFFSR_165 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_1_BUFX2_95 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_1_NAND3X1_56 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_2_OAI22X1_38 AND2X2_38/B DFFSR_23/S FILL
XFILL_45_DFFSR_196 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_45_1_0 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_0_NAND3X1_59 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_8_DFFSR_272 INVX1_3/gnd DFFSR_23/S FILL
XFILL_1_OAI22X1_41 INVX1_39/gnd DFFSR_54/S FILL
XFILL_35_DFFSR_199 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_0_OAI21X1_105 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_23_DFFPOSX1_35 INVX1_39/gnd DFFSR_54/S FILL
XFILL_0_OAI22X1_44 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_25_DFFSR_202 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_43_3_1 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_49_DFFSR_77 BUFX2_98/A DFFSR_32/S FILL
XFILL_7_8 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_7_NAND3X1_238 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_15_DFFSR_205 INVX1_3/gnd DFFSR_79/S FILL
XFILL_41_5_2 BUFX2_98/A DFFSR_32/S FILL
XINVX1_61 INVX1_61/A INVX1_39/gnd INVX1_61/Y DFFSR_54/S INVX1
XFILL_33_DFFSR_27 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_5_DFFSR_74 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_22_DFFSR_67 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_48_DFFSR_123 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_38_DFFSR_126 BUFX2_99/A DFFSR_7/S FILL
XINVX1_179 INVX1_179/A DFFSR_8/gnd INVX1_179/Y DFFSR_8/S INVX1
XFILL_8_NAND3X1_172 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_4_BUFX2_12 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_1_DFFSR_202 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_28_DFFSR_129 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_9_XOR2X1_4 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_42_DFFSR_233 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_1_NAND2X1_153 BUFX2_98/A DFFSR_32/S FILL
XFILL_4_INVX1_176 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_4_DFFSR_4 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_18_DFFSR_132 INVX1_3/gnd DFFSR_79/S FILL
XFILL_32_DFFSR_236 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_22_DFFSR_239 INVX1_39/gnd DFFSR_54/S FILL
XFILL_4_NAND3X1_11 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_9_NAND3X1_106 INVX1_3/gnd DFFSR_23/S FILL
XFILL_2_INVX1_68 INVX1_67/gnd DFFSR_201/S FILL
XFILL_30_DFFSR_74 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_3_XNOR2X1_2 BUFX2_98/A DFFSR_6/S FILL
XFILL_41_DFFSR_34 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_3_NOR2X1_11 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_13_DFFPOSX1_10 INVX1_67/gnd DFFSR_201/S FILL
XFILL_12_DFFSR_242 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_3_NAND3X1_14 DFFSR_4/gnd DFFSR_4/S FILL
XDFFSR_132 DFFSR_156/D CLKBUF1_18/Y BUFX2_61/Y DFFSR_79/S BUFX2_85/A INVX1_3/gnd DFFSR_79/S
+ DFFSR
XFILL_2_NAND3X1_17 BUFX2_99/A DFFSR_7/S FILL
XFILL_14_DFFSR_24 BUFX2_98/A DFFSR_6/S FILL
XFILL_4_DFFSR_129 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_2_OR2X2_4 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_1_BUFX2_59 AND2X2_38/B DFFSR_23/S FILL
XFILL_1_NAND3X1_20 BUFX2_99/A DFFSR_7/S FILL
XFILL_45_DFFSR_160 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_11_AOI22X1_7 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_0_NAND3X1_23 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_15_XOR2X1_11 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_8_DFFSR_236 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_35_DFFSR_163 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_5_NOR3X1_5 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_49_DFFSR_267 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_28_DFFSR_8 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_25_DFFSR_166 AND2X2_38/B DFFSR_59/S FILL
XFILL_49_DFFSR_41 BUFX2_98/A DFFSR_6/S FILL
XFILL_1_INVX1_213 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_38_DFFSR_81 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_39_DFFSR_270 INVX1_39/gnd DFFSR_54/S FILL
XFILL_51_0_2 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_7_NAND3X1_202 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_15_DFFSR_169 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_7_AOI22X1_1 INVX1_1/gnd DFFSR_97/S FILL
XFILL_29_DFFSR_273 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_3_DFFPOSX1_21 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_19_DFFSR_276 BUFX2_72/gnd DFFSR_276/S FILL
XINVX1_25 INVX1_25/A DFFSR_8/gnd INVX1_25/Y DFFSR_60/S INVX1
XDFFSR_78 DFFSR_78/Q DFFSR_45/CLK DFFSR_15/R DFFSR_4/S DFFSR_70/Q OR2X2_3/gnd DFFSR_4/S
+ DFFSR
XFILL_5_DFFSR_38 BUFX2_98/A DFFSR_6/S FILL
XFILL_22_DFFSR_31 BUFX2_79/A DFFSR_6/S FILL
XFILL_11_DFFSR_71 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_0_NOR2X1_48 INVX1_39/gnd DFFSR_34/S FILL
XFILL_8_NAND3X1_136 DFFSR_1/gnd DFFSR_81/S FILL
XINVX1_143 INVX1_143/A BUFX2_8/gnd INVX1_143/Y DFFSR_81/S INVX1
XFILL_1_DFFSR_166 AND2X2_38/B DFFSR_59/S FILL
XFILL_12_DFFPOSX1_40 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_1_NAND2X1_117 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_42_DFFSR_197 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_15_XOR2X1_1 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_49_DFFSR_4 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_46_DFFSR_88 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_5_DFFSR_273 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_32_DFFSR_200 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_22_DFFSR_203 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_2_INVX1_32 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_2_DFFSR_85 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_19_DFFSR_78 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_30_DFFSR_38 BUFX2_98/A DFFSR_6/S FILL
XFILL_12_DFFSR_206 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_17_1_1 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_22_DFFPOSX1_29 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_15_CLKBUF1_1 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_1_BUFX2_23 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_6_NAND3X1_232 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_15_3_2 INVX1_39/gnd DFFSR_34/S FILL
XFILL_4_INVX1_6 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_45_DFFSR_124 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_8_DFFSR_200 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_35_DFFSR_127 BUFX2_99/A DFFSR_92/S FILL
XFILL_11_NOR3X1_2 INVX1_1/gnd DFFSR_53/S FILL
XFILL_49_DFFSR_231 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_25_DFFSR_130 BUFX2_79/A DFFSR_6/S FILL
XFILL_38_DFFSR_45 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_1_INVX1_177 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_39_DFFSR_234 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_27_DFFSR_85 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_15_DFFSR_133 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_7_NAND3X1_166 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_29_DFFSR_237 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_0_NAND2X1_147 OR2X2_2/gnd DFFSR_216/S FILL
XDFFSR_42 DFFSR_42/Q DFFSR_7/CLK DFFSR_9/R DFFSR_32/S DFFSR_34/Q OR2X2_4/gnd DFFSR_32/S
+ DFFSR
XFILL_19_DFFSR_240 INVX1_39/gnd DFFSR_34/S FILL
XFILL_11_DFFSR_35 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_0_XNOR2X1_3 INVX1_1/gnd DFFSR_97/S FILL
XFILL_0_NOR2X1_12 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_8_NAND3X1_100 AND2X2_38/B DFFSR_59/S FILL
XINVX1_107 DFFSR_207/Q DFFSR_34/gnd INVX1_107/Y DFFSR_34/S INVX1
XFILL_1_DFFSR_130 BUFX2_79/A DFFSR_6/S FILL
XFILL_15_DFFSR_2 BUFX2_79/A DFFSR_7/S FILL
XFILL_42_DFFSR_161 INVX1_67/gnd DFFSR_175/S FILL
XFILL_42_6_0 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_46_DFFSR_52 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_35_DFFSR_92 BUFX2_99/A DFFSR_92/S FILL
XFILL_5_DFFSR_237 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_12_XOR2X1_12 INVX1_3/gnd DFFSR_23/S FILL
XFILL_32_DFFSR_164 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_46_DFFSR_268 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_22_DFFSR_167 OR2X2_2/gnd DFFSR_216/S FILL
XAOI22X1_5 NOR3X1_2/Y AOI22X1_5/B DFFSR_93/Q NOR3X1_1/Y DFFSR_8/gnd AOI22X1_5/Y DFFSR_60/S
+ AOI22X1
XFILL_19_DFFSR_42 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_2_DFFSR_49 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_36_DFFSR_271 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_6_BUFX2_77 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_12_DFFSR_170 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_26_DFFSR_274 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_4_AOI22X1_2 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_8_OAI21X1_118 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_16_DFFSR_277 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_20_CLKBUF1_32 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_6_NAND3X1_196 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_2_DFFPOSX1_15 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_19_CLKBUF1_35 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_43_DFFSR_99 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_8_DFFSR_164 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_18_CLKBUF1_38 OR2X2_3/gnd DFFSR_60/S FILL
XAND2X2_11 AND2X2_11/A AND2X2_11/B BUFX2_99/A AND2X2_11/Y DFFSR_7/S AND2X2
XFILL_49_DFFSR_195 DFFSR_46/gnd DFFSR_62/S FILL
XNAND3X1_232 NAND3X1_228/Y NAND3X1_229/Y INVX1_178/Y DFFSR_4/gnd NAND3X1_236/B DFFSR_98/S
+ NAND3X1
XFILL_4_AND2X2_8 BUFX2_99/A DFFSR_7/S FILL
XFILL_1_INVX1_141 INVX1_67/gnd DFFSR_201/S FILL
XFILL_39_DFFSR_198 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_17_CLKBUF1_41 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_27_DFFSR_49 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_16_DFFSR_89 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_2_DFFSR_274 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_7_NAND3X1_130 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_29_DFFSR_201 INVX1_67/gnd DFFSR_201/S FILL
XFILL_16_CLKBUF1_44 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_11_DFFPOSX1_34 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_19_DFFSR_204 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_0_NAND2X1_111 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_15_CLKBUF1_47 BUFX2_98/A DFFSR_32/S FILL
XFILL_52_1_0 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_4_NOR2X1_83 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_12_CLKBUF1_2 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_42_DFFSR_125 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_21_DFFPOSX1_23 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_46_DFFSR_16 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_35_DFFSR_56 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_24_DFFSR_96 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_5_DFFSR_201 INVX1_67/gnd DFFSR_201/S FILL
XFILL_50_3_1 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_32_DFFSR_128 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_46_DFFSR_232 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_5_NAND3X1_226 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_22_DFFSR_131 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_36_DFFSR_235 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_2_DFFSR_13 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_1_DFFPOSX1_45 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_48_5_2 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_6_BUFX2_41 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_12_DFFSR_134 INVX1_1/gnd DFFSR_53/S FILL
XFILL_26_DFFSR_238 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_11_6 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_7_XNOR2X1_1 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_28_1 INVX1_3/gnd DFFSR_79/S FILL
XFILL_16_DFFSR_241 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_6_NAND3X1_160 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_43_DFFSR_63 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_4_INVX1_97 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_8_DFFSR_128 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_49_DFFSR_159 DFFSR_62/gnd DFFSR_208/S FILL
XNAND3X1_196 INVX1_163/A NAND2X1_91/Y OAI21X1_55/Y DFFSR_46/gnd NAND3X1_196/Y DFFSR_62/S
+ NAND3X1
XFILL_39_DFFSR_162 BUFX2_99/A DFFSR_92/S FILL
XFILL_1_INVX1_105 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_27_DFFSR_13 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_16_DFFSR_53 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_2_DFFSR_238 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_16_4_0 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_3_BUFX2_88 INVX1_3/gnd DFFSR_23/S FILL
XFILL_29_DFFSR_165 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_43_DFFSR_269 INVX1_67/gnd DFFSR_201/S FILL
XFILL_19_DFFSR_168 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_15_CLKBUF1_11 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_33_DFFSR_272 INVX1_3/gnd DFFSR_23/S FILL
XNOR2X1_50 NOR2X1_50/A NOR2X1_50/B INVX1_39/gnd NOR2X1_50/Y DFFSR_34/S NOR2X1
XFILL_14_6_1 INVX1_39/gnd DFFSR_54/S FILL
XFILL_14_CLKBUF1_14 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_3_DFFSR_1 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_23_DFFSR_275 BUFX2_99/A DFFSR_92/S FILL
XFILL_1_AOI22X1_3 INVX1_1/gnd DFFSR_97/S FILL
XFILL_4_NOR2X1_47 AND2X2_38/B DFFSR_23/S FILL
XFILL_13_CLKBUF1_17 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_13_DFFSR_278 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_12_CLKBUF1_20 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_7_OAI21X1_112 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_24_DFFSR_60 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_11_CLKBUF1_23 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_35_DFFSR_20 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_7_DFFSR_67 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_5_DFFSR_165 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_46_DFFSR_196 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_10_CLKBUF1_26 INVX1_1/gnd DFFSR_53/S FILL
XFILL_5_NAND3X1_190 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_9_DFFSR_272 INVX1_3/gnd DFFSR_23/S FILL
XFILL_1_OR2X2_1 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_36_DFFSR_199 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_9_CLKBUF1_29 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_26_DFFSR_202 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_16_DFFSR_205 INVX1_3/gnd DFFSR_79/S FILL
XFILL_27_DFFSR_5 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_8_CLKBUF1_32 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_6_NAND3X1_124 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_7_CLKBUF1_35 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_10_DFFPOSX1_28 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_43_DFFSR_27 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_4_INVX1_61 INVX1_39/gnd DFFSR_54/S FILL
XFILL_32_DFFSR_67 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_6_CLKBUF1_38 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_7_10 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_49_DFFSR_123 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_5_CLKBUF1_41 OR2X2_4/gnd DFFSR_3/S FILL
XNAND3X1_160 INVX1_151/A AOI22X1_21/C NAND2X1_74/Y OR2X2_1/gnd AOI21X1_10/A DFFSR_51/S
+ NAND3X1
XFILL_39_DFFSR_126 BUFX2_99/A DFFSR_7/S FILL
XCLKBUF1_38 BUFX2_1/Y OR2X2_3/gnd CLKBUF1_38/Y DFFSR_60/S CLKBUF1
XFILL_16_DFFSR_17 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_2_DFFSR_202 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_4_CLKBUF1_44 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_3_BUFX2_52 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_29_DFFSR_129 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_24_1_1 AND2X2_38/B DFFSR_59/S FILL
XFILL_43_DFFSR_233 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_3_CLKBUF1_47 BUFX2_98/A DFFSR_32/S FILL
XFILL_20_DFFPOSX1_17 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_19_DFFSR_132 INVX1_3/gnd DFFSR_79/S FILL
XFILL_6_0_0 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_33_DFFSR_236 DFFSR_62/gnd DFFSR_62/S FILL
XNOR2X1_14 NOR2X1_14/A NOR2X1_14/B INVX1_1/gnd NOR2X1_14/Y DFFSR_97/S NOR2X1
XFILL_48_DFFSR_1 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_22_3_2 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_23_DFFSR_239 INVX1_39/gnd DFFSR_54/S FILL
XFILL_4_NAND3X1_220 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_40_DFFSR_74 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_4_XNOR2X1_2 BUFX2_98/A DFFSR_6/S FILL
XFILL_4_NOR2X1_11 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_13_DFFSR_242 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_4_2_1 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_0_DFFPOSX1_39 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_50_1 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_24_DFFSR_24 BUFX2_98/A DFFSR_6/S FILL
XFILL_7_DFFSR_31 BUFX2_79/A DFFSR_6/S FILL
XFILL_5_DFFSR_129 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_13_DFFSR_64 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_2_4_2 INVX1_67/gnd DFFSR_201/S FILL
XFILL_0_BUFX2_99 BUFX2_99/A DFFSR_7/S FILL
XFILL_46_DFFSR_160 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_5_NAND3X1_154 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_9_DFFSR_236 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_36_DFFSR_163 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_3_INVX1_3 INVX1_3/gnd DFFSR_79/S FILL
XFILL_50_DFFSR_267 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_26_DFFSR_166 AND2X2_38/B DFFSR_59/S FILL
XFILL_0_XOR2X1_1 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_2_INVX1_213 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_48_DFFSR_81 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_40_DFFSR_270 INVX1_39/gnd DFFSR_54/S FILL
XFILL_16_DFFSR_169 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_8_AOI22X1_1 INVX1_1/gnd DFFSR_97/S FILL
XFILL_30_DFFSR_273 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_20_DFFSR_276 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_4_INVX1_25 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_4_DFFSR_78 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_49_6_0 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_32_DFFSR_31 BUFX2_79/A DFFSR_6/S FILL
XFILL_19_DFFPOSX1_47 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_21_DFFSR_71 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_1_NOR2X1_48 INVX1_39/gnd DFFSR_34/S FILL
XFILL_10_DFFSR_279 BUFX2_99/A DFFSR_7/S FILL
XNAND3X1_124 NAND2X1_52/Y NAND3X1_124/B AND2X2_26/Y XOR2X1_4/gnd NOR2X1_58/A DFFSR_97/S
+ NAND3X1
XFILL_2_DFFSR_166 AND2X2_38/B DFFSR_59/S FILL
XFILL_3_BUFX2_16 BUFX2_98/A DFFSR_32/S FILL
XFILL_8_XOR2X1_8 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_43_DFFSR_197 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_3_CLKBUF1_11 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_6_DFFSR_273 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_6_OAI21X1_106 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_2_CLKBUF1_14 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_33_DFFSR_200 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_4_NAND3X1_184 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_1_CLKBUF1_17 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_23_DFFSR_203 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_29_DFFSR_78 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_40_DFFSR_38 BUFX2_98/A DFFSR_6/S FILL
XFILL_1_INVX1_72 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_13_DFFSR_206 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_0_CLKBUF1_20 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_16_CLKBUF1_1 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_13_DFFSR_28 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_0_BUFX2_63 BUFX2_98/A DFFSR_32/S FILL
XFILL_46_DFFSR_124 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_5_NAND3X1_118 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_9_DFFSR_200 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_36_DFFSR_127 BUFX2_99/A DFFSR_92/S FILL
XFILL_50_DFFSR_231 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_26_DFFSR_130 BUFX2_79/A DFFSR_6/S FILL
XFILL_48_DFFSR_45 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_2_INVX1_177 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_40_DFFSR_234 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_37_DFFSR_85 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_16_DFFSR_133 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_30_DFFSR_237 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_20_DFFSR_240 INVX1_39/gnd DFFSR_34/S FILL
XFILL_4_DFFSR_42 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_21_DFFSR_35 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_19_DFFPOSX1_11 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_1_XNOR2X1_3 INVX1_1/gnd DFFSR_97/S FILL
XFILL_10_DFFSR_75 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_1_NOR2X1_12 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_10_DFFSR_243 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_3_NAND3X1_214 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_2_DFFSR_130 BUFX2_79/A DFFSR_6/S FILL
XFILL_43_DFFSR_161 INVX1_67/gnd DFFSR_175/S FILL
XFILL_14_XOR2X1_5 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_39_DFFSR_8 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_55_6 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_45_DFFSR_92 BUFX2_99/A DFFSR_92/S FILL
XFILL_26_DFFPOSX1_2 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_6_DFFSR_237 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_13_XOR2X1_12 INVX1_3/gnd DFFSR_23/S FILL
XFILL_33_DFFSR_164 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_47_DFFSR_268 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_25_DFFPOSX1_5 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_23_DFFSR_167 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_6_AND2X2_1 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_4_NAND3X1_148 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_1_INVX1_36 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_29_DFFSR_42 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_1_DFFSR_89 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_37_DFFSR_271 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_18_DFFSR_82 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_24_DFFPOSX1_8 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_13_DFFSR_170 OR2X2_6/gnd DFFSR_92/S FILL
XOAI21X1_106 DFFSR_208/S INVX1_204/Y OAI21X1_106/C XOR2X1_1/gnd DFFSR_278/D DFFSR_208/S
+ OAI21X1
XFILL_27_DFFSR_274 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_5_AOI22X1_2 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_9_DFFPOSX1_22 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_17_DFFSR_277 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_0_BUFX2_27 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_23_4_0 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_9_DFFSR_164 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_18_DFFPOSX1_41 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_10_NOR3X1_6 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_50_DFFSR_195 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_21_6_1 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_2_INVX1_141 INVX1_67/gnd DFFSR_201/S FILL
XFILL_40_DFFSR_198 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_9_DFFSR_96 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_37_DFFSR_49 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_26_DFFSR_89 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_2_NAND3X1_244 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_3_DFFSR_274 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_3_5_0 INVX1_67/gnd DFFSR_175/S FILL
XFILL_30_DFFSR_201 INVX1_67/gnd DFFSR_201/S FILL
XFILL_20_DFFSR_204 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_10_DFFSR_39 INVX1_3/gnd DFFSR_79/S FILL
XFILL_5_OAI21X1_100 INVX1_3/gnd DFFSR_79/S FILL
XFILL_10_DFFSR_207 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_5_NOR2X1_83 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_3_NAND3X1_178 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_13_CLKBUF1_2 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_43_DFFSR_125 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_45_DFFSR_56 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_34_DFFSR_96 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_6_DFFSR_201 INVX1_67/gnd DFFSR_201/S FILL
XFILL_33_DFFSR_128 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_47_DFFSR_232 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_23_DFFSR_131 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_4_NAND3X1_112 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_37_DFFSR_235 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_1_DFFSR_53 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_18_DFFSR_46 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_13_DFFSR_134 INVX1_1/gnd DFFSR_53/S FILL
XFILL_5_BUFX2_81 BUFX2_79/A DFFSR_7/S FILL
XFILL_15_3 INVX1_39/gnd DFFSR_54/S FILL
XFILL_27_DFFSR_238 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_6_NAND2X1_148 INVX1_67/gnd DFFSR_175/S FILL
XFILL_8_XNOR2X1_1 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_17_DFFSR_241 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_26_DFFSR_2 BUFX2_79/A DFFSR_7/S FILL
XFILL_31_1_1 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_9_DFFSR_128 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_50_DFFSR_159 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_2_INVX1_105 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_9_DFFSR_60 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_40_DFFSR_162 BUFX2_99/A DFFSR_92/S FILL
XFILL_15_DFFSR_93 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_37_DFFSR_13 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_26_DFFSR_53 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_29_3_2 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_3_DFFSR_238 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_2_NAND3X1_208 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_10_XOR2X1_13 INVX1_1/gnd DFFSR_97/S FILL
XFILL_30_DFFSR_165 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_44_DFFSR_269 INVX1_67/gnd DFFSR_201/S FILL
XFILL_20_DFFSR_168 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_34_DFFSR_272 INVX1_3/gnd DFFSR_23/S FILL
XFILL_10_DFFSR_171 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_24_DFFSR_275 BUFX2_99/A DFFSR_92/S FILL
XFILL_2_AOI22X1_3 INVX1_1/gnd DFFSR_97/S FILL
XFILL_9_4_2 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_3_NAND3X1_142 INVX1_67/gnd DFFSR_175/S FILL
XFILL_5_NOR2X1_47 AND2X2_38/B DFFSR_23/S FILL
XFILL_14_DFFSR_278 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_14_DFFPOSX1_2 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_8_DFFPOSX1_16 INVX1_67/gnd DFFSR_175/S FILL
XFILL_13_DFFPOSX1_5 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_34_DFFSR_60 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_45_DFFSR_20 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_5_NAND2X1_178 INVX1_1/gnd DFFSR_53/S FILL
XFILL_6_DFFSR_165 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_12_DFFPOSX1_8 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_47_DFFSR_196 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_1_DFFSR_17 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_37_DFFSR_199 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_18_DFFSR_10 DFFSR_5/gnd DFFSR_5/S FILL
XBUFX2_85 BUFX2_85/A XOR2X1_4/gnd BUFX2_85/Y DFFSR_97/S BUFX2
XFILL_5_BUFX2_45 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_0_DFFSR_275 BUFX2_99/A DFFSR_92/S FILL
XFILL_27_DFFSR_202 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_17_DFFPOSX1_35 INVX1_39/gnd DFFSR_54/S FILL
XFILL_6_NAND2X1_112 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_17_DFFSR_205 INVX1_3/gnd DFFSR_79/S FILL
XFILL_1_NAND3X1_238 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_9_AOI21X1_37 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_42_DFFSR_67 DFFSR_34/gnd DFFSR_34/S FILL
XNAND2X1_148 DFFPOSX1_28/Q INVX1_208/Y INVX1_67/gnd AOI21X1_50/A DFFSR_175/S NAND2X1
XFILL_10_CLKBUF1_3 BUFX2_98/A DFFSR_6/S FILL
XFILL_50_DFFSR_123 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_8_AOI21X1_40 INVX1_39/gnd DFFSR_54/S FILL
XFILL_27_DFFPOSX1_24 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_9_DFFSR_24 BUFX2_98/A DFFSR_6/S FILL
XFILL_40_DFFSR_126 BUFX2_99/A DFFSR_7/S FILL
XFILL_26_DFFSR_17 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_15_DFFSR_57 BUFX2_79/A DFFSR_6/S FILL
XFILL_7_AOI21X1_43 INVX1_3/gnd DFFSR_79/S FILL
XFILL_3_DFFSR_202 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_2_NAND3X1_172 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_2_BUFX2_92 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_30_DFFSR_129 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_6_AOI21X1_46 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_44_DFFSR_233 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_20_DFFSR_132 INVX1_3/gnd DFFSR_79/S FILL
XFILL_7_DFFPOSX1_46 INVX1_39/gnd DFFSR_34/S FILL
XFILL_5_AOI21X1_49 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_34_DFFSR_236 DFFSR_62/gnd DFFSR_62/S FILL
XAOI21X1_46 AOI21X1_46/A AOI21X1_46/B BUFX2_39/Y BUFX2_7/gnd AOI21X1_46/Y DFFSR_151/S
+ AOI21X1
XFILL_10_DFFSR_135 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_4_AOI21X1_52 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_24_DFFSR_239 INVX1_39/gnd DFFSR_54/S FILL
XFILL_50_DFFSR_74 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_5_XNOR2X1_2 BUFX2_98/A DFFSR_6/S FILL
XFILL_5_NOR2X1_11 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_3_NAND3X1_106 INVX1_3/gnd DFFSR_23/S FILL
XFILL_3_AOI21X1_55 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_14_DFFSR_242 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_37_3 BUFX2_99/A DFFSR_92/S FILL
XFILL_2_AOI21X1_58 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_5_NAND2X1_142 INVX1_67/gnd DFFSR_175/S FILL
XFILL_34_DFFSR_24 BUFX2_98/A DFFSR_6/S FILL
XFILL_6_DFFSR_71 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_6_DFFSR_129 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_23_DFFSR_64 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_1_AOI21X1_61 AND2X2_38/B DFFSR_59/S FILL
XFILL_47_DFFSR_160 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_0_AOI21X1_64 AND2X2_38/B DFFSR_59/S FILL
XFILL_37_DFFSR_163 DFFSR_1/gnd DFFSR_1/S FILL
XBUFX2_49 INVX1_59/Y INVX1_1/gnd BUFX2_49/Y DFFSR_97/S BUFX2
XFILL_0_DFFSR_239 INVX1_39/gnd DFFSR_54/S FILL
XFILL_27_DFFSR_166 AND2X2_38/B DFFSR_59/S FILL
XFILL_3_INVX1_213 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_41_DFFSR_270 INVX1_39/gnd DFFSR_54/S FILL
XFILL_17_DFFSR_169 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_17_DFFSR_9 BUFX2_79/A DFFSR_6/S FILL
XFILL_8_OAI21X1_88 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_9_AOI22X1_1 INVX1_1/gnd DFFSR_97/S FILL
XFILL_31_DFFSR_273 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_1_NAND3X1_202 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_21_DFFSR_276 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_7_OAI21X1_91 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_3_INVX1_65 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_42_DFFSR_31 BUFX2_79/A DFFSR_6/S FILL
XFILL_31_DFFSR_71 XOR2X1_4/gnd DFFSR_91/S FILL
XNAND2X1_112 OR2X2_4/B OR2X2_4/A OR2X2_4/gnd AOI21X1_44/B DFFSR_3/S NAND2X1
XFILL_2_NOR2X1_48 INVX1_39/gnd DFFSR_34/S FILL
XFILL_6_OAI21X1_94 INVX1_67/gnd DFFSR_175/S FILL
XFILL_11_DFFSR_279 BUFX2_99/A DFFSR_7/S FILL
XFILL_5_OAI21X1_97 BUFX2_72/gnd DFFSR_276/S FILL
XOAI21X1_94 BUFX2_54/Y INVX1_191/Y OAI21X1_94/C INVX1_67/gnd DFFSR_266/D DFFSR_175/S
+ OAI21X1
XFILL_15_DFFSR_21 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_3_DFFSR_166 AND2X2_38/B DFFSR_59/S FILL
XFILL_2_NAND3X1_136 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_2_BUFX2_56 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_6_AOI21X1_10 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_44_DFFSR_197 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_7_DFFPOSX1_10 INVX1_67/gnd DFFSR_201/S FILL
XFILL_5_AOI21X1_13 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_7_DFFSR_273 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_6_NOR3X1_2 INVX1_1/gnd DFFSR_53/S FILL
XFILL_4_NAND2X1_172 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_34_DFFSR_200 DFFSR_62/gnd DFFSR_62/S FILL
XAOI21X1_10 AOI21X1_10/A AOI21X1_10/B AOI21X1_10/C BUFX2_8/gnd OAI21X1_41/B DFFSR_81/S
+ AOI21X1
XFILL_38_DFFSR_5 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_4_AOI21X1_16 INVX1_67/gnd DFFSR_175/S FILL
XFILL_24_DFFSR_203 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_39_DFFSR_78 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_50_DFFSR_38 BUFX2_98/A DFFSR_6/S FILL
XFILL_30_4_0 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_2_DFFPOSX1_2 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_3_AOI21X1_19 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_14_DFFSR_206 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_16_DFFPOSX1_29 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_1_DFFPOSX1_5 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_2_AOI21X1_22 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_17_CLKBUF1_1 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_6_DFFSR_35 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_5_NAND2X1_106 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_28_6_1 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_23_DFFSR_28 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_0_DFFPOSX1_8 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_12_DFFSR_68 BUFX2_98/A DFFSR_6/S FILL
XFILL_1_AOI21X1_25 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_0_NAND3X1_232 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_47_DFFSR_124 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_0_AOI21X1_28 AND2X2_38/B DFFSR_23/S FILL
XFILL_37_DFFSR_127 BUFX2_99/A DFFSR_92/S FILL
XBUFX2_13 AND2X2_1/Y DFFSR_28/gnd BUFX2_13/Y DFFSR_8/S BUFX2
XFILL_0_DFFSR_203 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_27_DFFSR_130 BUFX2_79/A DFFSR_6/S FILL
XFILL_3_INVX1_177 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_41_DFFSR_234 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_26_DFFPOSX1_18 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_47_DFFSR_85 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_17_DFFSR_133 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_31_DFFSR_237 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_1_NAND3X1_166 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_8_OAI21X1_52 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_6_NAND2X1_73 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_21_DFFSR_240 INVX1_39/gnd DFFSR_34/S FILL
XFILL_7_OAI21X1_55 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_31_DFFSR_35 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_3_INVX1_29 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_3_DFFSR_82 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_2_XNOR2X1_3 INVX1_1/gnd DFFSR_97/S FILL
XFILL_20_DFFSR_75 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_2_NOR2X1_12 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_6_DFFPOSX1_40 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_5_NAND2X1_76 INVX1_3/gnd DFFSR_23/S FILL
XFILL_6_OAI21X1_58 INVX1_39/gnd DFFSR_54/S FILL
XFILL_11_DFFSR_243 BUFX2_7/gnd DFFSR_151/S FILL
XNAND2X1_73 INVX1_145/A INVX1_175/A OR2X2_1/gnd INVX1_151/A DFFSR_59/S NAND2X1
XFILL_5_OAI21X1_61 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_4_NAND2X1_79 XOR2X1_1/gnd DFFSR_151/S FILL
XOAI21X1_58 OAI21X1_73/A OAI21X1_73/B OAI21X1_58/C INVX1_39/gnd AOI21X1_29/A DFFSR_54/S
+ OAI21X1
XFILL_3_DFFSR_130 BUFX2_79/A DFFSR_6/S FILL
XFILL_2_NAND3X1_100 AND2X2_38/B DFFSR_59/S FILL
XFILL_2_BUFX2_20 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_4_OAI21X1_64 INVX1_1/gnd DFFSR_53/S FILL
XFILL_3_NAND2X1_82 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_44_DFFSR_161 INVX1_67/gnd DFFSR_175/S FILL
XFILL_10_AOI22X1_8 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_3_OAI21X1_67 INVX1_1/gnd DFFSR_97/S FILL
XFILL_2_NAND2X1_85 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_7_DFFSR_237 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_14_XOR2X1_12 INVX1_3/gnd DFFSR_23/S FILL
XFILL_4_NAND2X1_136 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_34_DFFSR_164 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_2_OAI21X1_70 INVX1_3/gnd DFFSR_23/S FILL
XFILL_1_NAND2X1_88 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_48_DFFSR_268 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_24_DFFSR_167 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_0_NAND2X1_91 INVX1_39/gnd DFFSR_54/S FILL
XFILL_39_DFFSR_42 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_0_INVX1_214 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_38_DFFSR_271 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_0_INVX1_76 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_1_OAI21X1_73 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_28_DFFSR_82 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_14_DFFSR_170 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_38_1_1 BUFX2_79/A DFFSR_7/S FILL
XFILL_28_DFFSR_274 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_6_AOI22X1_2 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_0_OAI21X1_76 INVX1_1/gnd DFFSR_53/S FILL
XFILL_2_OAI21X1_118 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_25_DFFPOSX1_48 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_18_DFFSR_277 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_12_DFFSR_32 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_36_3_2 BUFX2_99/A DFFSR_92/S FILL
XFILL_0_NAND3X1_196 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_5_DFFSR_8 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_0_DFFSR_167 OR2X2_2/gnd DFFSR_216/S FILL
XDFFSR_277 BUFX2_75/A CLKBUF1_15/Y DFFSR_274/R DFFSR_201/S DFFSR_277/D BUFX2_72/gnd
+ DFFSR_201/S DFFSR
XFILL_3_INVX1_141 INVX1_67/gnd DFFSR_201/S FILL
XFILL_41_DFFSR_198 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_47_DFFSR_49 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_36_DFFSR_89 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_4_DFFSR_274 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_31_DFFSR_201 INVX1_67/gnd DFFSR_201/S FILL
XFILL_8_OAI21X1_16 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_1_NAND3X1_130 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_6_NAND2X1_37 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_21_DFFSR_204 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_7_OAI21X1_19 BUFX2_98/A DFFSR_32/S FILL
XFILL_20_DFFSR_39 INVX1_3/gnd DFFSR_79/S FILL
XFILL_3_DFFSR_46 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_5_NAND2X1_40 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_3_NAND2X1_166 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_6_OAI21X1_22 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_11_DFFSR_207 DFFSR_62/gnd DFFSR_62/S FILL
XNAND2X1_37 DFFSR_161/Q AND2X2_18/Y BUFX2_7/gnd NAND2X1_37/Y DFFSR_216/S NAND2X1
XFILL_4_NAND2X1_43 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_5_OAI21X1_25 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_6_NOR2X1_83 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_14_CLKBUF1_2 BUFX2_72/gnd DFFSR_276/S FILL
XOAI21X1_22 XOR2X1_1/B NOR2X1_66/B OAI21X1_22/C DFFSR_34/gnd XOR2X1_2/A DFFSR_34/S
+ OAI21X1
XFILL_4_OAI21X1_28 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_3_NAND2X1_46 INVX1_39/gnd DFFSR_34/S FILL
XDFFPOSX1_40 INVX1_175/A CLKBUF1_48/Y NOR2X1_76/Y OR2X2_1/gnd DFFSR_59/S DFFPOSX1
XFILL_44_DFFSR_125 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_13_XOR2X1_9 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_15_DFFPOSX1_23 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_2_NAND2X1_49 INVX1_3/gnd DFFSR_79/S FILL
XFILL_3_OAI21X1_31 AND2X2_38/B DFFSR_23/S FILL
XFILL_7_DFFSR_201 INVX1_67/gnd DFFSR_201/S FILL
XFILL_44_DFFSR_96 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_34_DFFSR_128 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_4_NAND2X1_100 INVX1_39/gnd DFFSR_54/S FILL
XFILL_2_OAI21X1_34 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_1_NAND2X1_52 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_48_DFFSR_232 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_24_DFFSR_131 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_5_AND2X2_5 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_1_OAI21X1_37 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_0_NAND2X1_55 INVX1_39/gnd DFFSR_34/S FILL
XFILL_38_DFFSR_235 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_0_DFFSR_93 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_0_INVX1_40 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_0_INVX1_178 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_17_DFFSR_86 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_28_DFFSR_46 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_14_DFFSR_134 INVX1_1/gnd DFFSR_53/S FILL
XFILL_28_DFFSR_238 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_0_OAI21X1_40 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_9_XNOR2X1_1 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_25_DFFPOSX1_12 AND2X2_38/B DFFSR_23/S FILL
XFILL_18_DFFSR_241 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_0_NAND3X1_160 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_50_DFFSR_8 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_7_AOI22X1_12 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_5_DFFPOSX1_34 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_0_DFFSR_131 NOR3X1_6/gnd DFFSR_79/S FILL
XDFFSR_241 INVX1_68/A CLKBUF1_2/Y BUFX2_67/Y DFFSR_201/S DFFSR_241/D BUFX2_72/gnd
+ DFFSR_201/S DFFSR
XFILL_6_AOI22X1_15 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_3_INVX1_105 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_41_DFFSR_162 BUFX2_99/A DFFSR_92/S FILL
XFILL_25_DFFSR_93 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_47_DFFSR_13 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_36_DFFSR_53 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_5_AOI22X1_18 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_4_DFFSR_238 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_11_XOR2X1_13 INVX1_1/gnd DFFSR_97/S FILL
XFILL_31_DFFSR_165 BUFX2_72/gnd DFFSR_201/S FILL
XAOI22X1_15 NOR3X1_4/Y DFFSR_231/Q DFFSR_231/D NOR3X1_3/Y DFFSR_46/gnd AOI22X1_15/Y
+ DFFSR_54/S AOI22X1
XFILL_45_DFFSR_269 INVX1_67/gnd DFFSR_201/S FILL
XFILL_4_AOI22X1_21 AND2X2_38/B DFFSR_59/S FILL
XFILL_21_DFFSR_168 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_3_DFFSR_10 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_35_DFFSR_272 INVX1_3/gnd DFFSR_23/S FILL
XFILL_3_AOI22X1_24 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_3_NAND2X1_130 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_11_DFFSR_171 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_25_DFFSR_275 BUFX2_99/A DFFSR_92/S FILL
XFILL_2_AOI22X1_27 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_3_AOI22X1_3 INVX1_1/gnd DFFSR_97/S FILL
XFILL_6_NOR2X1_47 AND2X2_38/B DFFSR_23/S FILL
XFILL_15_DFFSR_278 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_3_NAND2X1_10 BUFX2_79/A DFFSR_7/S FILL
XFILL_10_OAI22X1_51 INVX1_39/gnd DFFSR_54/S FILL
XFILL_2_NAND2X1_13 BUFX2_99/A DFFSR_92/S FILL
XFILL_10_1_2 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_7_DFFSR_165 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_44_DFFSR_60 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_1_OAI21X1_112 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_24_DFFPOSX1_42 INVX1_39/gnd DFFSR_34/S FILL
XFILL_1_NAND2X1_16 BUFX2_79/A DFFSR_7/S FILL
XFILL_48_DFFSR_196 XOR2X1_1/gnd DFFSR_151/S FILL
XAND2X2_9 AND2X2_9/A AND2X2_9/B DFFSR_28/gnd AND2X2_9/Y DFFSR_3/S AND2X2
XFILL_8_NAND3X1_72 INVX1_39/gnd DFFSR_34/S FILL
XFILL_0_NAND2X1_19 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_8_NAND3X1_245 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_0_DFFSR_57 BUFX2_79/A DFFSR_6/S FILL
XFILL_0_INVX1_142 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_38_DFFSR_199 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_28_DFFSR_10 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_17_DFFSR_50 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_7_NAND3X1_75 BUFX2_79/A DFFSR_7/S FILL
XFILL_1_DFFSR_275 BUFX2_99/A DFFSR_92/S FILL
XFILL_4_BUFX2_85 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_28_DFFSR_202 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_6_NAND3X1_78 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_18_DFFSR_205 INVX1_3/gnd DFFSR_79/S FILL
XFILL_5_NAND3X1_81 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_0_NAND3X1_124 XOR2X1_4/gnd DFFSR_97/S FILL
XNAND3X1_78 DFFSR_194/Q BUFX2_30/Y NOR2X1_31/Y NOR3X1_6/gnd NAND3X1_78/Y DFFSR_79/S
+ NAND3X1
XFILL_16_DFFSR_6 BUFX2_79/A DFFSR_6/S FILL
XFILL_4_NAND3X1_84 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_11_CLKBUF1_3 BUFX2_98/A DFFSR_6/S FILL
XFILL_51_DFFSR_123 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_3_NAND3X1_87 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_2_NAND2X1_160 NOR3X1_6/gnd DFFSR_79/S FILL
XDFFSR_205 INVX1_93/A CLKBUF1_22/Y BUFX2_61/Y DFFSR_79/S DFFSR_205/D INVX1_3/gnd DFFSR_79/S
+ DFFSR
XFILL_41_DFFSR_126 BUFX2_99/A DFFSR_7/S FILL
XFILL_2_NAND3X1_90 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_36_DFFSR_17 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_8_DFFSR_64 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_25_DFFSR_57 BUFX2_79/A DFFSR_6/S FILL
XFILL_14_DFFSR_97 INVX1_1/gnd DFFSR_97/S FILL
XFILL_37_4_0 BUFX2_99/A DFFSR_7/S FILL
XFILL_4_DFFSR_202 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_31_DFFSR_129 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_1_NAND3X1_93 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_45_DFFSR_233 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_0_BUFX2_7 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_21_DFFSR_132 INVX1_3/gnd DFFSR_79/S FILL
XFILL_0_NAND3X1_96 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_14_DFFPOSX1_17 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_35_DFFSR_236 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_35_6_1 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_11_DFFSR_135 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_25_DFFSR_239 INVX1_39/gnd DFFSR_54/S FILL
XFILL_6_XNOR2X1_2 BUFX2_98/A DFFSR_6/S FILL
XFILL_6_NOR2X1_11 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_24_5 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_11_OAI22X1_12 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_15_DFFSR_242 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_37_DFFSR_2 BUFX2_79/A DFFSR_7/S FILL
XFILL_10_OAI22X1_15 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_44_DFFSR_24 BUFX2_98/A DFFSR_6/S FILL
XINVX1_98 INVX1_98/A DFFSR_46/gnd INVX1_98/Y DFFSR_62/S INVX1
XFILL_7_DFFSR_129 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_33_DFFSR_64 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_9_NAND3X1_33 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_48_DFFSR_160 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_9_OAI22X1_18 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_8_NAND3X1_36 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_0_INVX1_106 INVX1_67/gnd DFFSR_201/S FILL
XFILL_0_DFFSR_21 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_38_DFFSR_163 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_8_NAND3X1_209 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_17_DFFSR_14 INVX1_1/gnd DFFSR_53/S FILL
XINVX1_216 XOR2X1_13/A INVX1_1/gnd NOR2X1_81/A DFFSR_97/S INVX1
XFILL_7_NAND3X1_39 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_8_OAI22X1_21 BUFX2_98/A DFFSR_32/S FILL
XFILL_4_BUFX2_49 INVX1_1/gnd DFFSR_97/S FILL
XFILL_1_DFFSR_239 INVX1_39/gnd DFFSR_54/S FILL
XFILL_4_DFFPOSX1_28 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_28_DFFSR_166 AND2X2_38/B DFFSR_59/S FILL
XFILL_4_INVX1_213 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_42_DFFSR_270 INVX1_39/gnd DFFSR_54/S FILL
XFILL_7_OAI22X1_24 BUFX2_98/A DFFSR_32/S FILL
XFILL_6_NAND3X1_42 BUFX2_79/A DFFSR_6/S FILL
XFILL_18_DFFSR_169 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_32_DFFSR_273 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_6_OAI22X1_27 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_5_NAND3X1_45 OR2X2_3/gnd DFFSR_60/S FILL
XXOR2X1_11 XOR2X1_11/A INVX1_215/A XOR2X1_4/gnd XOR2X1_12/B DFFSR_91/S XOR2X1
XNAND3X1_42 DFFSR_6/Q NOR2X1_4/Y BUFX2_18/Y BUFX2_79/A AND2X2_11/B DFFSR_6/S NAND3X1
XFILL_22_DFFSR_276 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_4_NAND3X1_48 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_0_AOI22X1_4 BUFX2_99/A DFFSR_92/S FILL
XFILL_5_OAI22X1_30 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_41_DFFSR_71 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_3_NOR2X1_48 INVX1_39/gnd DFFSR_34/S FILL
XOAI22X1_27 INVX1_66/Y OAI22X1_45/B INVX1_67/Y OAI22X1_45/D OR2X2_2/gnd NOR2X1_35/A
+ DFFSR_216/S OAI22X1
XFILL_13_DFFPOSX1_47 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_12_DFFSR_279 BUFX2_99/A DFFSR_7/S FILL
XFILL_3_NAND3X1_51 BUFX2_99/A DFFSR_7/S FILL
XFILL_4_OAI22X1_33 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_2_NAND2X1_124 OR2X2_2/gnd DFFSR_216/S FILL
XDFFSR_169 DFFSR_169/Q CLKBUF1_11/Y BUFX2_69/Y DFFSR_62/S DFFSR_161/Q DFFSR_62/gnd
+ DFFSR_62/S DFFSR
XFILL_3_OAI22X1_36 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_2_NAND3X1_54 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_8_DFFSR_28 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_25_DFFSR_21 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_14_DFFSR_61 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_4_DFFSR_166 AND2X2_38/B DFFSR_59/S FILL
XFILL_1_NAND3X1_57 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_2_OAI22X1_39 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_1_BUFX2_96 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_45_1_1 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_45_DFFSR_197 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_0_NAND3X1_60 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_1_OAI22X1_42 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_8_DFFSR_273 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_35_DFFSR_200 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_0_AND2X2_10 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_0_OAI21X1_106 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_23_DFFPOSX1_36 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_0_OAI22X1_45 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_25_DFFSR_203 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_43_3_2 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_49_DFFSR_78 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_15_DFFSR_206 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_7_9 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_7_NAND3X1_239 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_18_CLKBUF1_1 DFFSR_8/gnd DFFSR_8/S FILL
XINVX1_62 INVX1_62/A DFFSR_62/gnd NOR3X1_3/B DFFSR_62/S INVX1
XFILL_33_DFFSR_28 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_22_DFFSR_68 BUFX2_98/A DFFSR_6/S FILL
XFILL_5_DFFSR_75 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_48_DFFSR_124 OR2X2_1/gnd DFFSR_59/S FILL
XINVX1_180 INVX1_180/A BUFX2_98/A INVX1_180/Y DFFSR_6/S INVX1
XFILL_38_DFFSR_127 BUFX2_99/A DFFSR_92/S FILL
XFILL_8_NAND3X1_173 XOR2X1_4/gnd DFFSR_91/S FILL
XCLKBUF1_1 BUFX2_2/Y DFFSR_8/gnd DFFSR_3/CLK DFFSR_8/S CLKBUF1
XFILL_4_BUFX2_13 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_1_DFFSR_203 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_28_DFFSR_130 BUFX2_79/A DFFSR_6/S FILL
XFILL_9_XOR2X1_5 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_1_NAND2X1_154 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_42_DFFSR_234 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_11_2_0 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_4_DFFSR_5 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_18_DFFSR_133 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_32_DFFSR_237 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_4_NAND3X1_12 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_22_DFFSR_240 INVX1_39/gnd DFFSR_34/S FILL
XFILL_41_DFFSR_35 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_3_XNOR2X1_3 INVX1_1/gnd DFFSR_97/S FILL
XFILL_2_INVX1_69 INVX1_3/gnd DFFSR_23/S FILL
XFILL_3_NOR2X1_12 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_30_DFFSR_75 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_13_DFFPOSX1_11 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_12_DFFSR_243 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_3_NAND3X1_15 DFFSR_4/gnd DFFSR_4/S FILL
XDFFSR_133 DFFSR_157/D DFFSR_5/CLK BUFX2_65/Y DFFSR_5/S BUFX2_86/A BUFX2_77/gnd DFFSR_5/S
+ DFFSR
XFILL_2_NAND3X1_18 BUFX2_79/A DFFSR_7/S FILL
XFILL_14_DFFSR_25 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_4_DFFSR_130 BUFX2_79/A DFFSR_6/S FILL
XFILL_1_BUFX2_60 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_1_NAND3X1_21 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_2_OR2X2_5 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_45_DFFSR_161 INVX1_67/gnd DFFSR_175/S FILL
XFILL_0_NAND3X1_24 INVX1_1/gnd DFFSR_97/S FILL
XFILL_15_XOR2X1_12 INVX1_3/gnd DFFSR_23/S FILL
XFILL_8_DFFSR_237 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_35_DFFSR_164 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_5_NOR3X1_6 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_49_DFFSR_268 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_28_DFFSR_9 BUFX2_79/A DFFSR_6/S FILL
XFILL_25_DFFSR_167 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_39_DFFSR_271 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_38_DFFSR_82 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_49_DFFSR_42 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_1_INVX1_214 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_15_DFFSR_170 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_7_NAND3X1_203 INVX1_1/gnd DFFSR_97/S FILL
XFILL_29_DFFSR_274 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_7_AOI22X1_2 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_3_DFFPOSX1_22 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_19_DFFSR_277 BUFX2_72/gnd DFFSR_201/S FILL
XINVX1_26 INVX1_26/A OR2X2_6/gnd INVX1_26/Y DFFSR_92/S INVX1
XDFFSR_79 DFFSR_79/Q DFFSR_79/CLK DFFSR_7/R DFFSR_79/S DFFSR_79/D NOR3X1_6/gnd DFFSR_79/S
+ DFFSR
XFILL_5_DFFSR_39 INVX1_3/gnd DFFSR_79/S FILL
XFILL_11_DFFSR_72 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_22_DFFSR_32 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_0_NOR2X1_49 AND2X2_38/B DFFSR_59/S FILL
XFILL_8_NAND3X1_137 BUFX2_7/gnd DFFSR_216/S FILL
XINVX1_144 INVX1_144/A BUFX2_8/gnd INVX1_144/Y DFFSR_51/S INVX1
XFILL_1_DFFSR_167 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_12_DFFPOSX1_41 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_15_XOR2X1_2 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_42_DFFSR_198 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_49_DFFSR_5 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_1_NAND2X1_118 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_46_DFFSR_89 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_5_DFFSR_274 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_32_DFFSR_201 INVX1_67/gnd DFFSR_201/S FILL
XFILL_22_DFFSR_204 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_2_INVX1_33 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_2_DFFSR_86 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_30_DFFSR_39 INVX1_3/gnd DFFSR_79/S FILL
XFILL_19_DFFSR_79 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_17_1_2 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_12_DFFSR_207 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_22_DFFPOSX1_30 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_15_CLKBUF1_2 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_1_BUFX2_24 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_6_NAND3X1_233 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_4_INVX1_7 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_45_DFFSR_125 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_8_DFFSR_201 INVX1_67/gnd DFFSR_201/S FILL
XFILL_35_DFFSR_128 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_11_NOR3X1_3 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_49_DFFSR_232 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_25_DFFSR_131 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_39_DFFSR_235 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_27_DFFSR_86 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_1_INVX1_178 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_38_DFFSR_46 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_15_DFFSR_134 INVX1_1/gnd DFFSR_53/S FILL
XFILL_7_NAND3X1_167 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_29_DFFSR_238 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_0_NAND2X1_148 INVX1_67/gnd DFFSR_175/S FILL
XFILL_19_DFFSR_241 BUFX2_72/gnd DFFSR_201/S FILL
XDFFSR_43 DFFSR_59/D DFFSR_57/CLK DFFSR_9/R DFFSR_6/S DFFSR_43/D BUFX2_98/A DFFSR_6/S
+ DFFSR
XFILL_11_DFFSR_36 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_0_XNOR2X1_4 BUFX2_98/A DFFSR_6/S FILL
XFILL_0_NOR2X1_13 BUFX2_99/A DFFSR_92/S FILL
XFILL_44_4_0 DFFSR_28/gnd DFFSR_3/S FILL
XINVX1_108 DFFSR_167/D BUFX2_77/gnd INVX1_108/Y DFFSR_5/S INVX1
XFILL_8_NAND3X1_101 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_1_DFFSR_131 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_15_DFFSR_3 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_42_6_1 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_4_INVX1_105 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_42_DFFSR_162 BUFX2_99/A DFFSR_92/S FILL
XFILL_46_DFFSR_53 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_35_DFFSR_93 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_5_DFFSR_238 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_12_XOR2X1_13 INVX1_1/gnd DFFSR_97/S FILL
XFILL_32_DFFSR_165 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_46_DFFSR_269 INVX1_67/gnd DFFSR_201/S FILL
XFILL_22_DFFSR_168 OR2X2_6/gnd DFFSR_92/S FILL
XAOI22X1_6 NOR3X1_2/Y DFFSR_110/D DFFSR_94/Q NOR3X1_1/Y DFFSR_4/gnd AOI22X1_6/Y DFFSR_4/S
+ AOI22X1
XFILL_2_DFFSR_50 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_36_DFFSR_272 INVX1_3/gnd DFFSR_23/S FILL
XFILL_19_DFFSR_43 BUFX2_98/A DFFSR_6/S FILL
XFILL_6_BUFX2_78 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_12_DFFSR_171 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_26_DFFSR_275 BUFX2_99/A DFFSR_92/S FILL
XFILL_4_AOI22X1_3 INVX1_1/gnd DFFSR_97/S FILL
XFILL_8_OAI21X1_119 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_16_DFFSR_278 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_20_CLKBUF1_33 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_6_NAND3X1_197 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_2_DFFPOSX1_16 INVX1_67/gnd DFFSR_175/S FILL
XFILL_19_CLKBUF1_36 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_8_DFFSR_165 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_49_DFFSR_196 XOR2X1_1/gnd DFFSR_151/S FILL
XAND2X2_12 AND2X2_12/A AND2X2_12/B BUFX2_98/A AND2X2_12/Y DFFSR_32/S AND2X2
XFILL_18_CLKBUF1_39 INVX1_1/gnd DFFSR_53/S FILL
XFILL_4_AND2X2_9 DFFSR_28/gnd DFFSR_3/S FILL
XNAND3X1_233 XOR2X1_7/Y NAND3X1_227/A NAND3X1_226/Y DFFSR_4/gnd NAND3X1_233/Y DFFSR_4/S
+ NAND3X1
XFILL_17_CLKBUF1_42 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_39_DFFSR_199 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_38_DFFSR_10 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_27_DFFSR_50 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_16_DFFSR_90 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_1_INVX1_142 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_6_1 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_2_DFFSR_275 BUFX2_99/A DFFSR_92/S FILL
XFILL_7_NAND3X1_131 AND2X2_38/B DFFSR_59/S FILL
XFILL_16_CLKBUF1_45 BUFX2_79/A DFFSR_7/S FILL
XFILL_29_DFFSR_202 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_11_DFFPOSX1_35 INVX1_39/gnd DFFSR_54/S FILL
XFILL_0_NAND2X1_112 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_15_CLKBUF1_48 INVX1_3/gnd DFFSR_79/S FILL
XFILL_19_DFFSR_205 INVX1_3/gnd DFFSR_79/S FILL
XFILL_52_1_1 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_12_CLKBUF1_3 BUFX2_98/A DFFSR_6/S FILL
XFILL_21_DFFPOSX1_24 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_42_DFFSR_126 BUFX2_99/A DFFSR_7/S FILL
XFILL_46_DFFSR_17 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_50_3_2 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_35_DFFSR_57 BUFX2_79/A DFFSR_6/S FILL
XFILL_24_DFFSR_97 INVX1_1/gnd DFFSR_97/S FILL
XFILL_5_DFFSR_202 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_32_DFFSR_129 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_46_DFFSR_233 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_5_NAND3X1_227 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_22_DFFSR_132 INVX1_3/gnd DFFSR_79/S FILL
XFILL_2_DFFSR_14 INVX1_1/gnd DFFSR_53/S FILL
XFILL_36_DFFSR_236 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_1_DFFPOSX1_46 INVX1_39/gnd DFFSR_34/S FILL
XFILL_6_BUFX2_42 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_12_DFFSR_135 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_26_DFFSR_239 INVX1_39/gnd DFFSR_54/S FILL
XFILL_11_7 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_7_XNOR2X1_2 BUFX2_98/A DFFSR_6/S FILL
XFILL_28_2 INVX1_3/gnd DFFSR_79/S FILL
XFILL_16_DFFSR_242 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_6_NAND3X1_161 AND2X2_38/B DFFSR_23/S FILL
XFILL_8_DFFSR_129 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_43_DFFSR_64 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_18_2_0 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_49_DFFSR_160 XOR2X1_4/gnd DFFSR_97/S FILL
XNAND3X1_197 INVX1_131/Y NAND3X1_196/Y OAI21X1_56/Y DFFSR_46/gnd OAI21X1_57/C DFFSR_54/S
+ NAND3X1
XFILL_1_INVX1_106 INVX1_67/gnd DFFSR_201/S FILL
XFILL_39_DFFSR_163 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_27_DFFSR_14 INVX1_1/gnd DFFSR_53/S FILL
XFILL_16_DFFSR_54 INVX1_39/gnd DFFSR_54/S FILL
XFILL_16_4_1 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_2_DFFSR_239 INVX1_39/gnd DFFSR_54/S FILL
XFILL_3_BUFX2_89 INVX1_1/gnd DFFSR_97/S FILL
XFILL_29_DFFSR_166 AND2X2_38/B DFFSR_59/S FILL
XFILL_43_DFFSR_270 INVX1_39/gnd DFFSR_54/S FILL
XFILL_15_CLKBUF1_12 AND2X2_38/B DFFSR_23/S FILL
XFILL_19_DFFSR_169 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_33_DFFSR_273 DFFSR_62/gnd DFFSR_208/S FILL
XNOR2X1_51 NOR2X1_51/A NOR2X1_51/B DFFSR_34/gnd NOR2X1_51/Y DFFSR_34/S NOR2X1
XFILL_14_6_2 INVX1_39/gnd DFFSR_54/S FILL
XFILL_14_CLKBUF1_15 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_3_DFFSR_2 BUFX2_79/A DFFSR_7/S FILL
XFILL_23_DFFSR_276 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_1_AOI22X1_4 BUFX2_99/A DFFSR_92/S FILL
XFILL_13_CLKBUF1_18 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_4_NOR2X1_48 INVX1_39/gnd DFFSR_34/S FILL
XFILL_13_DFFSR_279 BUFX2_99/A DFFSR_7/S FILL
XFILL_12_CLKBUF1_21 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_7_OAI21X1_113 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_7_DFFSR_68 BUFX2_98/A DFFSR_6/S FILL
XFILL_24_DFFSR_61 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_11_CLKBUF1_24 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_35_DFFSR_21 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_5_DFFSR_166 AND2X2_38/B DFFSR_59/S FILL
XFILL_5_NAND3X1_191 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_10_CLKBUF1_27 INVX1_1/gnd DFFSR_97/S FILL
XFILL_46_DFFSR_197 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_9_DFFSR_273 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_1_DFFPOSX1_10 INVX1_67/gnd DFFSR_201/S FILL
XFILL_36_DFFSR_200 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_1_OR2X2_2 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_1_AND2X2_10 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_9_CLKBUF1_30 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_26_DFFSR_203 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_16_DFFSR_206 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_8_CLKBUF1_33 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_27_DFFSR_6 BUFX2_79/A DFFSR_6/S FILL
XFILL_6_NAND3X1_125 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_7_CLKBUF1_36 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_10_DFFPOSX1_29 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_19_CLKBUF1_1 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_43_DFFSR_28 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_32_DFFSR_68 BUFX2_98/A DFFSR_6/S FILL
XFILL_6_CLKBUF1_39 INVX1_1/gnd DFFSR_53/S FILL
XFILL_49_DFFSR_124 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_5_CLKBUF1_42 DFFSR_4/gnd DFFSR_98/S FILL
XNAND3X1_161 INVX1_151/Y NAND3X1_158/B NAND2X1_78/Y AND2X2_38/B AOI21X1_10/B DFFSR_23/S
+ NAND3X1
XFILL_39_DFFSR_127 BUFX2_99/A DFFSR_92/S FILL
XCLKBUF1_39 BUFX2_6/Y INVX1_1/gnd CLKBUF1_39/Y DFFSR_53/S CLKBUF1
XFILL_16_DFFSR_18 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_4_CLKBUF1_45 BUFX2_79/A DFFSR_7/S FILL
XFILL_2_DFFSR_203 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_3_BUFX2_53 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_29_DFFSR_130 BUFX2_79/A DFFSR_6/S FILL
XFILL_24_1_2 AND2X2_38/B DFFSR_59/S FILL
XFILL_43_DFFSR_234 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_3_CLKBUF1_48 INVX1_3/gnd DFFSR_79/S FILL
XFILL_20_DFFPOSX1_18 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_19_DFFSR_133 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_33_DFFSR_237 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_6_0_1 BUFX2_7/gnd DFFSR_216/S FILL
XNOR2X1_15 NOR2X1_15/A NOR2X1_15/B BUFX2_99/A NOR2X1_15/Y DFFSR_7/S NOR2X1
XFILL_48_DFFSR_2 BUFX2_79/A DFFSR_7/S FILL
XFILL_23_DFFSR_240 INVX1_39/gnd DFFSR_34/S FILL
XFILL_4_NAND3X1_221 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_4_XNOR2X1_3 INVX1_1/gnd DFFSR_97/S FILL
XFILL_4_NOR2X1_12 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_40_DFFSR_75 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_13_DFFSR_243 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_0_DFFPOSX1_40 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_4_2_2 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_50_2 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_7_DFFSR_32 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_24_DFFSR_25 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_13_DFFSR_65 BUFX2_79/A DFFSR_7/S FILL
XFILL_5_DFFSR_130 BUFX2_79/A DFFSR_6/S FILL
XFILL_46_DFFSR_161 INVX1_67/gnd DFFSR_175/S FILL
XFILL_5_NAND3X1_155 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_9_DFFSR_237 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_36_DFFSR_164 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_3_INVX1_4 BUFX2_99/A DFFSR_7/S FILL
XFILL_50_DFFSR_268 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_26_DFFSR_167 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_0_XOR2X1_2 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_40_DFFSR_271 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_51_4_0 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_48_DFFSR_82 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_2_INVX1_214 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_16_DFFSR_170 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_30_DFFSR_274 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_8_AOI22X1_2 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_20_DFFSR_277 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_49_6_1 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_32_DFFSR_32 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_4_DFFSR_79 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_21_DFFSR_72 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_19_DFFPOSX1_48 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_1_NOR2X1_49 AND2X2_38/B DFFSR_59/S FILL
XFILL_10_DFFSR_280 OR2X2_6/gnd DFFSR_53/S FILL
XNAND3X1_125 DFFSR_200/D BUFX2_31/Y BUFX2_24/Y BUFX2_77/gnd NAND3X1_127/A DFFSR_98/S
+ NAND3X1
XFILL_2_DFFSR_167 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_3_BUFX2_17 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_8_XOR2X1_9 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_43_DFFSR_198 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_3_CLKBUF1_12 AND2X2_38/B DFFSR_23/S FILL
XFILL_6_DFFSR_274 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_6_OAI21X1_107 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_33_DFFSR_201 INVX1_67/gnd DFFSR_201/S FILL
XFILL_2_CLKBUF1_15 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_23_DFFSR_204 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_4_NAND3X1_185 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_1_CLKBUF1_18 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_29_DFFSR_79 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_40_DFFSR_39 INVX1_3/gnd DFFSR_79/S FILL
XFILL_1_INVX1_73 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_0_CLKBUF1_21 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_13_DFFSR_207 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_16_CLKBUF1_2 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_13_DFFSR_29 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_0_BUFX2_64 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_46_DFFSR_125 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_5_NAND3X1_119 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_9_DFFSR_201 INVX1_67/gnd DFFSR_201/S FILL
XFILL_36_DFFSR_128 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_50_DFFSR_232 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_26_DFFSR_131 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_40_DFFSR_235 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_37_DFFSR_86 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_2_INVX1_178 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_48_DFFSR_46 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_16_DFFSR_134 INVX1_1/gnd DFFSR_53/S FILL
XFILL_30_DFFSR_238 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_20_DFFSR_241 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_21_DFFSR_36 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_4_DFFSR_43 BUFX2_98/A DFFSR_6/S FILL
XFILL_1_XNOR2X1_4 BUFX2_98/A DFFSR_6/S FILL
XFILL_10_DFFSR_76 BUFX2_79/A DFFSR_7/S FILL
XFILL_19_DFFPOSX1_12 AND2X2_38/B DFFSR_23/S FILL
XFILL_1_NOR2X1_13 BUFX2_99/A DFFSR_92/S FILL
XFILL_10_DFFSR_244 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_3_NAND3X1_215 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_2_DFFSR_131 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_14_XOR2X1_6 BUFX2_99/A DFFSR_7/S FILL
XFILL_43_DFFSR_162 BUFX2_99/A DFFSR_92/S FILL
XFILL_55_7 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_39_DFFSR_9 BUFX2_79/A DFFSR_6/S FILL
XFILL_45_DFFSR_93 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_6_DFFSR_238 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_13_XOR2X1_13 INVX1_1/gnd DFFSR_97/S FILL
XFILL_26_DFFPOSX1_3 INVX1_39/gnd DFFSR_34/S FILL
XFILL_33_DFFSR_165 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_47_DFFSR_269 INVX1_67/gnd DFFSR_201/S FILL
XFILL_25_DFFPOSX1_6 AND2X2_38/B DFFSR_23/S FILL
XFILL_6_AND2X2_2 BUFX2_99/A DFFSR_7/S FILL
XFILL_23_DFFSR_168 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_4_NAND3X1_149 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_1_DFFSR_90 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_1_INVX1_37 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_29_DFFSR_43 BUFX2_98/A DFFSR_6/S FILL
XFILL_18_DFFSR_83 INVX1_3/gnd DFFSR_79/S FILL
XFILL_37_DFFSR_272 INVX1_3/gnd DFFSR_23/S FILL
XFILL_24_DFFPOSX1_9 INVX1_67/gnd DFFSR_201/S FILL
XFILL_13_DFFSR_171 BUFX2_8/gnd DFFSR_81/S FILL
XOAI21X1_107 DFFSR_91/S INVX1_205/Y OAI21X1_107/C OR2X2_6/gnd DFFSR_279/D DFFSR_92/S
+ OAI21X1
XFILL_25_2_0 AND2X2_38/B DFFSR_23/S FILL
XFILL_27_DFFSR_275 BUFX2_99/A DFFSR_92/S FILL
XFILL_5_AOI22X1_3 INVX1_1/gnd DFFSR_97/S FILL
XFILL_9_DFFPOSX1_23 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_17_DFFSR_278 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_0_BUFX2_28 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_23_4_1 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_9_DFFSR_165 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_5_3_0 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_18_DFFPOSX1_42 INVX1_39/gnd DFFSR_34/S FILL
XFILL_50_DFFSR_196 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_21_6_2 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_40_DFFSR_199 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_48_DFFSR_10 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_37_DFFSR_50 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_9_DFFSR_97 INVX1_1/gnd DFFSR_97/S FILL
XFILL_2_INVX1_142 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_26_DFFSR_90 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_2_NAND3X1_245 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_3_DFFSR_275 BUFX2_99/A DFFSR_92/S FILL
XFILL_3_5_1 INVX1_67/gnd DFFSR_175/S FILL
XFILL_30_DFFSR_202 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_20_DFFSR_205 INVX1_3/gnd DFFSR_79/S FILL
XFILL_10_DFFSR_40 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_5_OAI21X1_101 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_10_DFFSR_208 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_3_NAND3X1_179 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_13_CLKBUF1_3 BUFX2_98/A DFFSR_6/S FILL
XFILL_43_DFFSR_126 BUFX2_99/A DFFSR_7/S FILL
XFILL_45_DFFSR_57 BUFX2_79/A DFFSR_6/S FILL
XFILL_34_DFFSR_97 INVX1_1/gnd DFFSR_97/S FILL
XFILL_6_DFFSR_202 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_33_DFFSR_129 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_47_DFFSR_233 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_23_DFFSR_132 INVX1_3/gnd DFFSR_79/S FILL
XFILL_4_NAND3X1_113 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_37_DFFSR_236 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_18_DFFSR_47 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_1_DFFSR_54 INVX1_39/gnd DFFSR_54/S FILL
XFILL_5_BUFX2_82 INVX1_1/gnd DFFSR_97/S FILL
XFILL_13_DFFSR_135 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_15_4 INVX1_39/gnd DFFSR_54/S FILL
XFILL_27_DFFSR_239 INVX1_39/gnd DFFSR_54/S FILL
XFILL_8_XNOR2X1_2 BUFX2_98/A DFFSR_6/S FILL
XFILL_6_NAND2X1_149 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_17_DFFSR_242 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_26_DFFSR_3 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_31_1_2 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_9_DFFSR_129 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_50_DFFSR_160 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_40_DFFSR_163 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_2_INVX1_106 INVX1_67/gnd DFFSR_201/S FILL
XFILL_9_DFFSR_61 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_37_DFFSR_14 INVX1_1/gnd DFFSR_53/S FILL
XFILL_15_DFFSR_94 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_26_DFFSR_54 INVX1_39/gnd DFFSR_54/S FILL
XFILL_2_NAND3X1_209 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_3_DFFSR_239 INVX1_39/gnd DFFSR_54/S FILL
XFILL_10_XOR2X1_14 INVX1_1/gnd DFFSR_53/S FILL
XFILL_30_DFFSR_166 AND2X2_38/B DFFSR_59/S FILL
XFILL_44_DFFSR_270 INVX1_39/gnd DFFSR_54/S FILL
XFILL_20_DFFSR_169 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_34_DFFSR_273 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_10_DFFSR_172 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_24_DFFSR_276 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_2_AOI22X1_4 BUFX2_99/A DFFSR_92/S FILL
XFILL_3_NAND3X1_143 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_5_NOR2X1_48 INVX1_39/gnd DFFSR_34/S FILL
XFILL_14_DFFSR_279 BUFX2_99/A DFFSR_7/S FILL
XFILL_14_DFFPOSX1_3 INVX1_39/gnd DFFSR_34/S FILL
XFILL_8_DFFPOSX1_17 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_13_DFFPOSX1_6 AND2X2_38/B DFFSR_23/S FILL
XFILL_34_DFFSR_61 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_45_DFFSR_21 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_5_NAND2X1_179 INVX1_1/gnd DFFSR_97/S FILL
XFILL_6_DFFSR_166 AND2X2_38/B DFFSR_59/S FILL
XFILL_12_DFFPOSX1_9 INVX1_67/gnd DFFSR_201/S FILL
XFILL_47_DFFSR_197 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_37_DFFSR_200 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_1_DFFSR_18 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_18_DFFSR_11 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_2_AND2X2_10 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_0_DFFSR_276 BUFX2_72/gnd DFFSR_276/S FILL
XBUFX2_86 BUFX2_86/A BUFX2_77/gnd BUFX2_86/Y DFFSR_98/S BUFX2
XFILL_5_BUFX2_46 BUFX2_98/A DFFSR_6/S FILL
XFILL_17_DFFPOSX1_36 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_27_DFFSR_203 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_6_NAND2X1_113 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_2_INVX1_1 INVX1_1/gnd DFFSR_53/S FILL
XFILL_17_DFFSR_206 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_1_NAND3X1_239 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_20_CLKBUF1_1 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_42_DFFSR_68 BUFX2_98/A DFFSR_6/S FILL
XNAND2X1_149 DFFSR_216/S NAND2X1_149/B OR2X2_2/gnd AOI21X1_50/B DFFSR_216/S NAND2X1
XFILL_10_CLKBUF1_4 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_50_DFFSR_124 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_8_AOI21X1_41 INVX1_39/gnd DFFSR_34/S FILL
XFILL_27_DFFPOSX1_25 BUFX2_79/A DFFSR_6/S FILL
XFILL_40_DFFSR_127 BUFX2_99/A DFFSR_92/S FILL
XFILL_7_AOI21X1_44 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_9_DFFSR_25 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_15_DFFSR_58 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_2_NAND3X1_173 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_26_DFFSR_18 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_3_DFFSR_203 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_30_DFFSR_130 BUFX2_79/A DFFSR_6/S FILL
XFILL_2_BUFX2_93 AND2X2_38/B DFFSR_59/S FILL
XFILL_6_AOI21X1_47 INVX1_67/gnd DFFSR_175/S FILL
XFILL_44_DFFSR_234 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_20_DFFSR_133 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_7_DFFPOSX1_47 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_5_AOI21X1_50 INVX1_67/gnd DFFSR_175/S FILL
XFILL_34_DFFSR_237 DFFSR_1/gnd DFFSR_1/S FILL
XAOI21X1_47 AOI21X1_47/A AOI21X1_47/B BUFX2_36/Y INVX1_67/gnd AOI21X1_47/Y DFFSR_175/S
+ AOI21X1
XFILL_10_DFFSR_136 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_4_AOI21X1_53 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_24_DFFSR_240 INVX1_39/gnd DFFSR_34/S FILL
XFILL_5_XNOR2X1_3 INVX1_1/gnd DFFSR_97/S FILL
XFILL_50_DFFSR_75 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_5_NOR2X1_12 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_3_AOI21X1_56 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_3_NAND3X1_107 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_14_DFFSR_243 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_37_4 BUFX2_99/A DFFSR_92/S FILL
XFILL_2_AOI21X1_59 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_5_NAND2X1_143 INVX1_67/gnd DFFSR_201/S FILL
XFILL_6_DFFSR_72 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_34_DFFSR_25 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_23_DFFSR_65 BUFX2_79/A DFFSR_7/S FILL
XFILL_6_DFFSR_130 BUFX2_79/A DFFSR_6/S FILL
XFILL_1_AOI21X1_62 INVX1_3/gnd DFFSR_23/S FILL
XFILL_47_DFFSR_161 INVX1_67/gnd DFFSR_175/S FILL
XFILL_0_AOI21X1_65 INVX1_3/gnd DFFSR_23/S FILL
XFILL_37_DFFSR_164 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_51_DFFSR_268 OR2X2_1/gnd DFFSR_51/S FILL
XBUFX2_50 INVX1_59/Y BUFX2_77/gnd DFFSR_8/R DFFSR_5/S BUFX2
XFILL_5_BUFX2_10 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_0_DFFSR_240 INVX1_39/gnd DFFSR_34/S FILL
XFILL_27_DFFSR_167 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_3_INVX1_214 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_41_DFFSR_271 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_17_DFFSR_170 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_8_OAI21X1_89 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_31_DFFSR_274 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_9_AOI22X1_2 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_1_NAND3X1_203 INVX1_1/gnd DFFSR_97/S FILL
XFILL_21_DFFSR_277 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_7_OAI21X1_92 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_3_INVX1_66 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_42_DFFSR_32 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_31_DFFSR_72 OR2X2_3/gnd DFFSR_60/S FILL
XNAND2X1_113 NAND3X1_245/Y NAND2X1_113/B OR2X2_4/gnd NAND2X1_113/Y DFFSR_3/S NAND2X1
XFILL_2_NOR2X1_49 AND2X2_38/B DFFSR_59/S FILL
XFILL_6_OAI21X1_95 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_11_DFFSR_280 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_5_OAI21X1_98 DFFSR_46/gnd DFFSR_54/S FILL
XOAI21X1_95 BUFX2_53/Y INVX1_192/Y OAI21X1_95/C BUFX2_7/gnd DFFSR_267/D DFFSR_216/S
+ OAI21X1
XFILL_2_NAND3X1_137 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_15_DFFSR_22 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_3_DFFSR_167 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_2_BUFX2_57 AND2X2_38/B DFFSR_23/S FILL
XFILL_44_DFFSR_198 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_6_AOI21X1_11 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_32_2_0 INVX1_1/gnd DFFSR_97/S FILL
XFILL_7_DFFSR_274 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_7_DFFPOSX1_11 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_4_NAND2X1_173 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_5_AOI21X1_14 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_34_DFFSR_201 INVX1_67/gnd DFFSR_201/S FILL
XFILL_6_NOR3X1_3 BUFX2_7/gnd DFFSR_216/S FILL
XAOI21X1_11 AOI21X1_11/A AOI21X1_11/B AOI21X1_11/C OR2X2_1/gnd OAI21X1_41/A DFFSR_51/S
+ AOI21X1
XFILL_38_DFFSR_6 BUFX2_79/A DFFSR_6/S FILL
XFILL_10_DFFSR_100 INVX1_1/gnd DFFSR_97/S FILL
XFILL_4_AOI21X1_17 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_24_DFFSR_204 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_30_4_1 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_39_DFFSR_79 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_50_DFFSR_39 INVX1_3/gnd DFFSR_79/S FILL
XFILL_3_AOI21X1_20 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_2_DFFPOSX1_3 INVX1_39/gnd DFFSR_34/S FILL
XFILL_14_DFFSR_207 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_1_DFFPOSX1_6 AND2X2_38/B DFFSR_23/S FILL
XFILL_16_DFFPOSX1_30 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_2_AOI21X1_23 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_17_CLKBUF1_2 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_5_NAND2X1_107 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_23_DFFSR_29 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_6_DFFSR_36 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_28_6_2 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_0_DFFPOSX1_9 INVX1_67/gnd DFFSR_201/S FILL
XFILL_12_DFFSR_69 BUFX2_98/A DFFSR_32/S FILL
XFILL_1_AOI21X1_26 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_0_NAND3X1_233 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_47_DFFSR_125 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_0_AOI21X1_29 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_37_DFFSR_128 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_51_DFFSR_232 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_0_DFFSR_204 BUFX2_7/gnd DFFSR_216/S FILL
XBUFX2_14 AND2X2_1/Y OR2X2_4/gnd BUFX2_14/Y DFFSR_32/S BUFX2
XFILL_27_DFFSR_131 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_41_DFFSR_235 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_26_DFFPOSX1_19 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_3_INVX1_178 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_47_DFFSR_86 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_17_DFFSR_134 INVX1_1/gnd DFFSR_53/S FILL
XFILL_8_OAI21X1_53 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_31_DFFSR_238 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_1_NAND3X1_167 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_6_NAND2X1_74 AND2X2_38/B DFFSR_59/S FILL
XFILL_7_OAI21X1_56 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_21_DFFSR_241 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_3_INVX1_30 INVX1_1/gnd DFFSR_53/S FILL
XFILL_3_DFFSR_83 INVX1_3/gnd DFFSR_79/S FILL
XFILL_31_DFFSR_36 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_2_XNOR2X1_4 BUFX2_98/A DFFSR_6/S FILL
XFILL_20_DFFSR_76 BUFX2_79/A DFFSR_7/S FILL
XFILL_6_DFFPOSX1_41 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_2_NOR2X1_13 BUFX2_99/A DFFSR_92/S FILL
XFILL_5_NAND2X1_77 AND2X2_38/B DFFSR_23/S FILL
XFILL_11_DFFSR_244 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_6_OAI21X1_59 DFFSR_62/gnd DFFSR_208/S FILL
XNAND2X1_74 AND2X2_32/Y AND2X2_33/Y AND2X2_38/B NAND2X1_74/Y DFFSR_59/S NAND2X1
XFILL_5_OAI21X1_62 INVX1_3/gnd DFFSR_79/S FILL
XFILL_4_NAND2X1_80 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_2_NAND3X1_101 XOR2X1_4/gnd DFFSR_91/S FILL
XOAI21X1_59 INVX1_157/A AOI21X1_29/Y OAI21X1_59/C DFFSR_62/gnd OAI21X1_59/Y DFFSR_208/S
+ OAI21X1
XFILL_4_OAI21X1_65 INVX1_1/gnd DFFSR_53/S FILL
XFILL_3_DFFSR_131 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_3_NAND2X1_83 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_2_BUFX2_21 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_44_DFFSR_162 BUFX2_99/A DFFSR_92/S FILL
XFILL_10_AOI22X1_9 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_2_NAND2X1_86 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_3_OAI21X1_68 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_7_DFFSR_238 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_14_XOR2X1_13 INVX1_1/gnd DFFSR_97/S FILL
XFILL_4_NAND2X1_137 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_34_DFFSR_165 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_48_DFFSR_269 INVX1_67/gnd DFFSR_201/S FILL
XFILL_2_OAI21X1_71 INVX1_3/gnd DFFSR_79/S FILL
XFILL_1_NAND2X1_89 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_24_DFFSR_168 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_0_NAND2X1_92 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_1_OAI21X1_74 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_39_DFFSR_43 BUFX2_98/A DFFSR_6/S FILL
XFILL_0_INVX1_215 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_28_DFFSR_83 INVX1_3/gnd DFFSR_79/S FILL
XFILL_38_DFFSR_272 INVX1_3/gnd DFFSR_23/S FILL
XFILL_0_INVX1_77 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_14_DFFSR_171 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_0_OAI21X1_77 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_38_1_2 BUFX2_79/A DFFSR_7/S FILL
XFILL_28_DFFSR_275 BUFX2_99/A DFFSR_92/S FILL
XFILL_6_AOI22X1_3 INVX1_1/gnd DFFSR_97/S FILL
XFILL_2_OAI21X1_119 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_25_DFFPOSX1_49 BUFX2_99/A DFFSR_92/S FILL
XFILL_18_DFFSR_278 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_12_DFFSR_33 BUFX2_98/A DFFSR_32/S FILL
XFILL_0_XOR2X1_10 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_0_NAND3X1_197 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_5_DFFSR_9 BUFX2_79/A DFFSR_6/S FILL
XFILL_51_DFFSR_196 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_0_DFFSR_168 OR2X2_6/gnd DFFSR_92/S FILL
XDFFSR_278 BUFX2_76/A CLKBUF1_15/Y DFFSR_274/R DFFSR_151/S DFFSR_278/D XOR2X1_1/gnd
+ DFFSR_151/S DFFSR
XFILL_41_DFFSR_199 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_47_DFFSR_50 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_3_INVX1_142 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_36_DFFSR_90 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_4_DFFSR_275 BUFX2_99/A DFFSR_92/S FILL
XFILL_8_OAI21X1_17 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_31_DFFSR_202 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_1_NAND3X1_131 AND2X2_38/B DFFSR_59/S FILL
XFILL_7_OAI21X1_20 AND2X2_38/B DFFSR_23/S FILL
XFILL_6_NAND2X1_38 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_21_DFFSR_205 INVX1_3/gnd DFFSR_79/S FILL
XFILL_3_DFFSR_47 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_20_DFFSR_40 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_6_OAI21X1_23 INVX1_67/gnd DFFSR_201/S FILL
XFILL_5_NAND2X1_41 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_3_NAND2X1_167 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_11_DFFSR_208 DFFSR_62/gnd DFFSR_208/S FILL
XNAND2X1_38 NOR3X1_4/A NOR3X1_4/B BUFX2_8/gnd NOR3X1_3/C DFFSR_81/S NAND2X1
XFILL_5_OAI21X1_26 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_4_NAND2X1_44 INVX1_39/gnd DFFSR_34/S FILL
XFILL_14_CLKBUF1_3 BUFX2_98/A DFFSR_6/S FILL
XOAI21X1_23 INVX1_131/Y XOR2X1_2/A OAI21X1_23/C INVX1_67/gnd OAI21X1_23/Y DFFSR_201/S
+ OAI21X1
XFILL_4_OAI21X1_29 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_3_NAND2X1_47 DFFSR_62/gnd DFFSR_208/S FILL
XDFFPOSX1_41 INVX1_159/A CLKBUF1_46/Y AOI21X1_63/Y DFFSR_8/gnd DFFSR_60/S DFFPOSX1
XFILL_44_DFFSR_126 BUFX2_99/A DFFSR_7/S FILL
XFILL_2_NAND2X1_50 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_44_DFFSR_97 INVX1_1/gnd DFFSR_97/S FILL
XFILL_3_OAI21X1_32 AND2X2_38/B DFFSR_59/S FILL
XFILL_15_DFFPOSX1_24 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_7_DFFSR_202 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_34_DFFSR_129 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_4_NAND2X1_101 INVX1_39/gnd DFFSR_54/S FILL
XFILL_48_DFFSR_233 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_2_OAI21X1_35 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_1_NAND2X1_53 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_5_AND2X2_6 BUFX2_99/A DFFSR_7/S FILL
XFILL_24_DFFSR_132 INVX1_3/gnd DFFSR_79/S FILL
XFILL_0_NAND2X1_56 AND2X2_38/B DFFSR_59/S FILL
XFILL_1_OAI21X1_38 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_0_INVX1_179 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_0_INVX1_41 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_28_DFFSR_47 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_0_DFFSR_94 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_38_DFFSR_236 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_17_DFFSR_87 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_19_1 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_14_DFFSR_135 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_0_OAI21X1_41 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_28_DFFSR_239 INVX1_39/gnd DFFSR_54/S FILL
XFILL_9_XNOR2X1_2 BUFX2_98/A DFFSR_6/S FILL
XFILL_18_DFFSR_242 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_25_DFFPOSX1_13 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_8_AOI22X1_10 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_0_NAND3X1_161 AND2X2_38/B DFFSR_23/S FILL
XFILL_50_DFFSR_9 BUFX2_79/A DFFSR_6/S FILL
XFILL_7_AOI22X1_13 AND2X2_38/B DFFSR_23/S FILL
XFILL_5_DFFPOSX1_35 INVX1_39/gnd DFFSR_54/S FILL
XDFFSR_242 INVX1_75/A DFFSR_5/CLK BUFX2_65/Y DFFSR_60/S DFFSR_242/D OR2X2_3/gnd DFFSR_60/S
+ DFFSR
XFILL_0_DFFSR_132 INVX1_3/gnd DFFSR_79/S FILL
XFILL_6_AOI22X1_16 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_41_DFFSR_163 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_3_INVX1_106 INVX1_67/gnd DFFSR_201/S FILL
XFILL_47_DFFSR_14 INVX1_1/gnd DFFSR_53/S FILL
XFILL_25_DFFSR_94 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_36_DFFSR_54 INVX1_39/gnd DFFSR_54/S FILL
XFILL_5_AOI22X1_19 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_4_DFFSR_239 INVX1_39/gnd DFFSR_54/S FILL
XFILL_11_XOR2X1_14 INVX1_1/gnd DFFSR_53/S FILL
XFILL_31_DFFSR_166 AND2X2_38/B DFFSR_59/S FILL
XAOI22X1_16 NOR3X1_4/Y DFFSR_232/Q DFFSR_224/Q NOR3X1_3/Y BUFX2_77/gnd AOI22X1_16/Y
+ DFFSR_5/S AOI22X1
XFILL_4_AOI22X1_22 INVX1_3/gnd DFFSR_79/S FILL
XFILL_45_DFFSR_270 INVX1_39/gnd DFFSR_54/S FILL
XFILL_21_DFFSR_169 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_3_DFFSR_11 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_35_DFFSR_273 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_3_AOI22X1_25 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_3_NAND2X1_131 INVX1_3/gnd DFFSR_79/S FILL
XFILL_11_DFFSR_172 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_25_DFFSR_276 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_3_AOI22X1_4 BUFX2_99/A DFFSR_92/S FILL
XFILL_2_AOI22X1_28 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_6_NOR2X1_48 INVX1_39/gnd DFFSR_34/S FILL
XFILL_15_DFFSR_279 BUFX2_99/A DFFSR_7/S FILL
XFILL_11_OAI22X1_49 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_3_NAND2X1_11 BUFX2_98/A DFFSR_6/S FILL
XFILL_10_OAI22X1_52 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_2_NAND2X1_14 BUFX2_98/A DFFSR_32/S FILL
XFILL_44_DFFSR_61 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_1_OAI21X1_113 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_7_DFFSR_166 AND2X2_38/B DFFSR_59/S FILL
XFILL_24_DFFPOSX1_43 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_9_NAND3X1_70 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_1_NAND2X1_17 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_48_DFFSR_197 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_8_NAND3X1_73 INVX1_1/gnd DFFSR_97/S FILL
XFILL_0_NAND2X1_20 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_8_NAND3X1_246 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_0_DFFSR_58 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_0_INVX1_143 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_28_DFFSR_11 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_38_DFFSR_200 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_3_AND2X2_10 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_17_DFFSR_51 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_1_DFFSR_276 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_7_NAND3X1_76 INVX1_1/gnd DFFSR_53/S FILL
XFILL_4_BUFX2_86 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_28_DFFSR_203 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_6_NAND3X1_79 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_18_DFFSR_206 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_5_NAND3X1_82 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_0_NAND3X1_125 BUFX2_77/gnd DFFSR_98/S FILL
XNAND3X1_79 NAND3X1_79/A NAND3X1_78/Y NAND3X1_79/C NOR3X1_6/gnd NOR2X1_40/B DFFSR_91/S
+ NAND3X1
XFILL_4_NAND3X1_85 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_16_DFFSR_7 BUFX2_79/A DFFSR_7/S FILL
XFILL_11_CLKBUF1_4 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_39_2_0 BUFX2_79/A DFFSR_6/S FILL
XFILL_3_NAND3X1_88 DFFSR_1/gnd DFFSR_81/S FILL
XDFFSR_206 DFFSR_214/D CLKBUF1_21/Y BUFX2_60/Y DFFSR_175/S DFFSR_206/D OR2X2_2/gnd
+ DFFSR_175/S DFFSR
XFILL_2_NAND2X1_161 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_41_DFFSR_127 BUFX2_99/A DFFSR_92/S FILL
XFILL_8_DFFSR_65 BUFX2_79/A DFFSR_7/S FILL
XFILL_2_NAND3X1_91 AND2X2_38/B DFFSR_59/S FILL
XFILL_25_DFFSR_58 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_14_DFFSR_98 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_36_DFFSR_18 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_4_DFFSR_203 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_37_4_1 BUFX2_99/A DFFSR_7/S FILL
XFILL_31_DFFSR_130 BUFX2_79/A DFFSR_6/S FILL
XFILL_1_NAND3X1_94 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_45_DFFSR_234 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_0_BUFX2_8 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_21_DFFSR_133 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_0_NAND3X1_97 AND2X2_38/B DFFSR_59/S FILL
XFILL_14_DFFPOSX1_18 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_35_DFFSR_237 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_35_6_2 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_11_DFFSR_136 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_25_DFFSR_240 INVX1_39/gnd DFFSR_34/S FILL
XFILL_6_XNOR2X1_3 INVX1_1/gnd DFFSR_97/S FILL
XFILL_6_NOR2X1_12 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_15_DFFSR_243 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_24_6 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_37_DFFSR_3 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_10_OAI22X1_16 AND2X2_38/B DFFSR_59/S FILL
XINVX1_99 INVX1_99/A DFFSR_46/gnd INVX1_99/Y DFFSR_62/S INVX1
XFILL_44_DFFSR_25 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_33_DFFSR_65 BUFX2_79/A DFFSR_7/S FILL
XFILL_7_DFFSR_130 BUFX2_79/A DFFSR_6/S FILL
XFILL_48_DFFSR_161 INVX1_67/gnd DFFSR_175/S FILL
XFILL_9_OAI22X1_19 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_8_NAND3X1_37 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_38_DFFSR_164 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_0_DFFSR_22 OR2X2_4/gnd DFFSR_32/S FILL
XINVX1_217 INVX1_217/A XOR2X1_4/gnd NOR2X1_81/B DFFSR_97/S INVX1
XFILL_8_NAND3X1_210 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_0_INVX1_107 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_17_DFFSR_15 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_8_OAI22X1_22 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_7_NAND3X1_40 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_1_DFFSR_240 INVX1_39/gnd DFFSR_34/S FILL
XFILL_4_BUFX2_50 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_4_DFFPOSX1_29 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_28_DFFSR_167 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_42_DFFSR_271 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_6_NAND3X1_43 BUFX2_99/A DFFSR_7/S FILL
XFILL_7_OAI22X1_25 INVX1_39/gnd DFFSR_54/S FILL
XFILL_18_DFFSR_170 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_32_DFFSR_274 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_5_NAND3X1_46 DFFSR_4/gnd DFFSR_4/S FILL
XXOR2X1_12 XOR2X1_12/A XOR2X1_12/B INVX1_3/gnd NOR2X1_79/B DFFSR_23/S XOR2X1
XFILL_6_OAI22X1_28 INVX1_3/gnd DFFSR_23/S FILL
XNAND3X1_43 BUFX2_87/A AND2X2_3/Y BUFX2_22/Y BUFX2_99/A AND2X2_11/A DFFSR_7/S NAND3X1
XFILL_22_DFFSR_277 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_0_AOI22X1_5 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_4_NAND3X1_49 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_5_OAI22X1_31 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_41_DFFSR_72 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_3_NOR2X1_49 AND2X2_38/B DFFSR_59/S FILL
XFILL_13_DFFPOSX1_48 XOR2X1_4/gnd DFFSR_97/S FILL
XOAI22X1_28 INVX1_69/Y OAI22X1_43/B INVX1_70/Y OAI22X1_43/D INVX1_3/gnd NOR2X1_38/B
+ DFFSR_23/S OAI22X1
XFILL_3_NAND3X1_52 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_12_DFFSR_280 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_4_OAI22X1_34 DFFSR_34/gnd DFFSR_1/S FILL
XDFFSR_170 DFFSR_170/Q CLKBUF1_3/Y BUFX2_63/Y DFFSR_92/S DFFSR_170/D OR2X2_6/gnd DFFSR_92/S
+ DFFSR
XFILL_2_NAND2X1_125 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_2_NAND3X1_55 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_8_DFFSR_29 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_3_OAI22X1_37 INVX1_3/gnd DFFSR_23/S FILL
XFILL_25_DFFSR_22 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_14_DFFSR_62 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_4_DFFSR_167 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_1_BUFX2_97 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_1_NAND3X1_58 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_2_OAI22X1_40 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_45_DFFSR_198 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_45_1_2 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_8_DFFSR_274 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_0_NAND3X1_61 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_1_OAI22X1_43 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_35_DFFSR_201 INVX1_67/gnd DFFSR_201/S FILL
XFILL_0_OAI21X1_107 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_0_AND2X2_11 BUFX2_99/A DFFSR_7/S FILL
XFILL_23_DFFPOSX1_37 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_11_DFFSR_100 INVX1_1/gnd DFFSR_97/S FILL
XFILL_0_OAI22X1_46 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_25_DFFSR_204 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_49_DFFSR_79 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_15_DFFSR_207 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_7_NAND3X1_240 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_18_CLKBUF1_2 BUFX2_72/gnd DFFSR_276/S FILL
XINVX1_63 NOR3X1_4/A XOR2X1_4/gnd INVX1_63/Y DFFSR_91/S INVX1
XFILL_33_DFFSR_29 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_5_DFFSR_76 BUFX2_79/A DFFSR_7/S FILL
XFILL_22_DFFSR_69 BUFX2_98/A DFFSR_32/S FILL
XFILL_48_DFFSR_125 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_13_0_0 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_38_DFFSR_128 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_8_NAND3X1_174 NOR3X1_6/gnd DFFSR_79/S FILL
XINVX1_181 DFFSR_1/D DFFSR_34/gnd INVX1_181/Y DFFSR_34/S INVX1
XCLKBUF1_2 BUFX2_5/Y BUFX2_72/gnd CLKBUF1_2/Y DFFSR_276/S CLKBUF1
XFILL_1_DFFSR_204 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_4_BUFX2_14 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_9_XOR2X1_6 BUFX2_99/A DFFSR_7/S FILL
XFILL_28_DFFSR_131 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_1_NAND2X1_155 BUFX2_79/A DFFSR_7/S FILL
XFILL_42_DFFSR_235 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_4_INVX1_178 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_11_2_1 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_4_DFFSR_6 BUFX2_79/A DFFSR_6/S FILL
XFILL_18_DFFSR_134 INVX1_1/gnd DFFSR_53/S FILL
XFILL_32_DFFSR_238 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_5_NAND3X1_10 BUFX2_79/A DFFSR_6/S FILL
XFILL_22_DFFSR_241 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_4_NAND3X1_13 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_9_NAND3X1_108 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_41_DFFSR_36 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_3_XNOR2X1_4 BUFX2_98/A DFFSR_6/S FILL
XFILL_30_DFFSR_76 BUFX2_79/A DFFSR_7/S FILL
XFILL_2_INVX1_70 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_3_NOR2X1_13 BUFX2_99/A DFFSR_92/S FILL
XFILL_13_DFFPOSX1_12 AND2X2_38/B DFFSR_23/S FILL
XFILL_12_DFFSR_244 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_3_NAND3X1_16 DFFSR_28/gnd DFFSR_8/S FILL
XDFFSR_134 DFFSR_158/D CLKBUF1_40/Y BUFX2_63/Y DFFSR_53/S BUFX2_87/A INVX1_1/gnd DFFSR_53/S
+ DFFSR
XFILL_2_NAND3X1_19 BUFX2_99/A DFFSR_92/S FILL
XFILL_14_DFFSR_26 BUFX2_79/A DFFSR_6/S FILL
XFILL_4_DFFSR_131 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_1_BUFX2_61 AND2X2_38/B DFFSR_59/S FILL
XFILL_2_OR2X2_6 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_1_NAND3X1_22 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_45_DFFSR_162 BUFX2_99/A DFFSR_92/S FILL
XFILL_11_AOI22X1_9 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_8_DFFSR_238 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_0_NAND3X1_25 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_15_XOR2X1_13 INVX1_1/gnd DFFSR_97/S FILL
XFILL_35_DFFSR_165 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_49_DFFSR_269 INVX1_67/gnd DFFSR_201/S FILL
XFILL_0_OAI22X1_10 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_25_DFFSR_168 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_49_DFFSR_43 BUFX2_98/A DFFSR_6/S FILL
XFILL_1_INVX1_215 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_39_DFFSR_272 INVX1_3/gnd DFFSR_23/S FILL
XFILL_38_DFFSR_83 INVX1_3/gnd DFFSR_79/S FILL
XFILL_15_DFFSR_171 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_7_NAND3X1_204 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_29_DFFSR_275 BUFX2_99/A DFFSR_92/S FILL
XFILL_7_AOI22X1_3 INVX1_1/gnd DFFSR_97/S FILL
XFILL_3_DFFPOSX1_23 NOR3X1_6/gnd DFFSR_91/S FILL
XDFFSR_80 DFFSR_80/Q DFFSR_45/CLK DFFSR_35/R DFFSR_4/S DFFSR_72/Q DFFSR_4/gnd DFFSR_4/S
+ DFFSR
XINVX1_27 DFFSR_84/D BUFX2_99/A INVX1_27/Y DFFSR_7/S INVX1
XFILL_19_DFFSR_278 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_5_DFFSR_40 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_22_DFFSR_33 BUFX2_98/A DFFSR_32/S FILL
XFILL_11_DFFSR_73 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_1_XOR2X1_10 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_0_NOR2X1_50 INVX1_39/gnd DFFSR_34/S FILL
XFILL_8_NAND3X1_138 INVX1_67/gnd DFFSR_201/S FILL
XINVX1_145 INVX1_145/A OR2X2_1/gnd INVX1_145/Y DFFSR_51/S INVX1
XFILL_1_DFFSR_168 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_12_DFFPOSX1_42 INVX1_39/gnd DFFSR_34/S FILL
XFILL_15_XOR2X1_3 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_1_NAND2X1_119 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_49_DFFSR_6 BUFX2_79/A DFFSR_6/S FILL
XFILL_4_INVX1_142 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_42_DFFSR_199 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_46_DFFSR_90 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_5_DFFSR_275 BUFX2_99/A DFFSR_92/S FILL
XFILL_32_DFFSR_202 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_22_DFFSR_205 INVX1_3/gnd DFFSR_79/S FILL
XFILL_30_DFFSR_40 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_19_DFFSR_80 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_2_DFFSR_87 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_2_INVX1_34 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_12_DFFSR_208 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_22_DFFPOSX1_31 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_15_CLKBUF1_3 BUFX2_98/A DFFSR_6/S FILL
XFILL_6_NAND3X1_234 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_1_BUFX2_25 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_4_INVX1_8 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_45_DFFSR_126 BUFX2_99/A DFFSR_7/S FILL
XFILL_8_DFFSR_202 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_35_DFFSR_129 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_11_NOR3X1_4 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_49_DFFSR_233 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_25_DFFSR_132 INVX1_3/gnd DFFSR_79/S FILL
XFILL_1_INVX1_179 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_38_DFFSR_47 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_39_DFFSR_236 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_27_DFFSR_87 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_15_DFFSR_135 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_7_NAND3X1_168 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_29_DFFSR_239 INVX1_39/gnd DFFSR_54/S FILL
XFILL_46_2_0 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_0_NAND2X1_149 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_19_DFFSR_242 OR2X2_3/gnd DFFSR_60/S FILL
XDFFSR_44 DFFSR_60/D CLKBUF1_37/Y DFFSR_8/R DFFSR_98/S DFFSR_44/D DFFSR_4/gnd DFFSR_98/S
+ DFFSR
XFILL_11_DFFSR_37 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_0_NOR2X1_14 INVX1_1/gnd DFFSR_97/S FILL
XFILL_44_4_1 DFFSR_28/gnd DFFSR_3/S FILL
XINVX1_109 DFFSR_151/D BUFX2_77/gnd INVX1_109/Y DFFSR_5/S INVX1
XFILL_8_NAND3X1_102 INVX1_3/gnd DFFSR_23/S FILL
XFILL_1_DFFSR_132 INVX1_3/gnd DFFSR_79/S FILL
XFILL_15_DFFSR_4 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_42_6_2 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_42_DFFSR_163 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_35_DFFSR_94 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_46_DFFSR_54 INVX1_39/gnd DFFSR_54/S FILL
XFILL_5_DFFSR_239 INVX1_39/gnd DFFSR_54/S FILL
XFILL_12_XOR2X1_14 INVX1_1/gnd DFFSR_53/S FILL
XFILL_32_DFFSR_166 AND2X2_38/B DFFSR_59/S FILL
XFILL_46_DFFSR_270 INVX1_39/gnd DFFSR_54/S FILL
XAOI22X1_7 NOR3X1_2/Y AOI22X1_7/B DFFSR_95/Q NOR3X1_1/Y DFFSR_8/gnd AOI22X1_7/Y DFFSR_8/S
+ AOI22X1
XFILL_22_DFFSR_169 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_19_DFFSR_44 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_2_DFFSR_51 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_36_DFFSR_273 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_12_DFFSR_172 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_6_BUFX2_79 BUFX2_79/A DFFSR_7/S FILL
XFILL_26_DFFSR_276 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_4_AOI22X1_4 BUFX2_99/A DFFSR_92/S FILL
XFILL_16_DFFSR_279 BUFX2_99/A DFFSR_7/S FILL
XFILL_20_CLKBUF1_34 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_6_NAND3X1_198 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_10_5_0 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_19_CLKBUF1_37 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_2_DFFPOSX1_17 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_8_DFFSR_166 AND2X2_38/B DFFSR_59/S FILL
XAND2X2_13 AND2X2_13/A AND2X2_13/B DFFSR_28/gnd AND2X2_13/Y DFFSR_3/S AND2X2
XFILL_49_DFFSR_197 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_18_CLKBUF1_40 OR2X2_6/gnd DFFSR_92/S FILL
XNAND3X1_234 NOR2X1_73/Y NAND3X1_233/Y NAND3X1_236/B BUFX2_77/gnd AOI21X1_36/B DFFSR_98/S
+ NAND3X1
XFILL_17_CLKBUF1_43 AND2X2_38/B DFFSR_23/S FILL
XFILL_1_INVX1_143 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_38_DFFSR_11 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_39_DFFSR_200 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_4_AND2X2_10 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_16_DFFSR_91 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_27_DFFSR_51 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_7_NAND3X1_132 AND2X2_38/B DFFSR_23/S FILL
XFILL_2_DFFSR_276 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_16_CLKBUF1_46 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_29_DFFSR_203 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_11_DFFPOSX1_36 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_19_DFFSR_206 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_0_NAND2X1_113 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_15_CLKBUF1_49 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_52_1_2 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_12_CLKBUF1_4 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_21_DFFPOSX1_25 BUFX2_79/A DFFSR_6/S FILL
XFILL_42_DFFSR_127 BUFX2_99/A DFFSR_92/S FILL
XFILL_35_DFFSR_58 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_46_DFFSR_18 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_24_DFFSR_98 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_5_DFFSR_203 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_32_DFFSR_130 BUFX2_79/A DFFSR_6/S FILL
XFILL_46_DFFSR_234 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_5_NAND3X1_228 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_22_DFFSR_133 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_2_DFFSR_15 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_1_DFFPOSX1_47 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_36_DFFSR_237 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_12_DFFSR_136 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_6_BUFX2_43 AND2X2_38/B DFFSR_23/S FILL
XFILL_26_DFFSR_240 INVX1_39/gnd DFFSR_34/S FILL
XFILL_7_XNOR2X1_3 INVX1_1/gnd DFFSR_97/S FILL
XFILL_16_DFFSR_243 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_20_0_0 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_6_NAND3X1_162 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_8_DFFSR_130 BUFX2_79/A DFFSR_6/S FILL
XFILL_43_DFFSR_65 BUFX2_79/A DFFSR_7/S FILL
XFILL_4_INVX1_99 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_18_2_1 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_49_DFFSR_161 INVX1_67/gnd DFFSR_175/S FILL
XFILL_0_1_0 BUFX2_72/gnd DFFSR_276/S FILL
XNAND3X1_198 AOI21X1_22/A AOI21X1_22/B AOI21X1_22/C DFFSR_62/gnd AOI21X1_29/B DFFSR_62/S
+ NAND3X1
XFILL_39_DFFSR_164 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_1_INVX1_107 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_27_DFFSR_15 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_16_DFFSR_55 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_16_4_2 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_3_BUFX2_90 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_2_DFFSR_240 INVX1_39/gnd DFFSR_34/S FILL
XFILL_16_CLKBUF1_10 INVX1_67/gnd DFFSR_201/S FILL
XFILL_29_DFFSR_167 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_43_DFFSR_271 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_15_CLKBUF1_13 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_19_DFFSR_170 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_33_DFFSR_274 BUFX2_72/gnd DFFSR_276/S FILL
XNOR2X1_52 NOR2X1_52/A NOR2X1_52/B DFFSR_1/gnd NOR2X1_52/Y DFFSR_1/S NOR2X1
XFILL_14_CLKBUF1_16 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_3_DFFSR_3 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_23_DFFSR_277 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_1_AOI22X1_5 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_51_DFFSR_72 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_4_NOR2X1_49 AND2X2_38/B DFFSR_59/S FILL
XFILL_13_CLKBUF1_19 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_13_DFFSR_280 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_12_CLKBUF1_22 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_7_OAI21X1_114 AND2X2_38/B DFFSR_59/S FILL
XFILL_11_CLKBUF1_25 INVX1_67/gnd DFFSR_201/S FILL
XFILL_35_DFFSR_22 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_7_DFFSR_69 BUFX2_98/A DFFSR_32/S FILL
XFILL_24_DFFSR_62 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_5_DFFSR_167 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_5_NAND3X1_192 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_46_DFFSR_198 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_10_CLKBUF1_28 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_9_DFFSR_274 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_36_DFFSR_201 INVX1_67/gnd DFFSR_201/S FILL
XFILL_1_OR2X2_3 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_1_DFFPOSX1_11 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_1_AND2X2_11 BUFX2_99/A DFFSR_7/S FILL
XFILL_12_DFFSR_100 INVX1_1/gnd DFFSR_97/S FILL
XFILL_26_DFFSR_204 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_9_CLKBUF1_31 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_16_DFFSR_207 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_8_CLKBUF1_34 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_27_DFFSR_7 BUFX2_79/A DFFSR_7/S FILL
XFILL_6_NAND3X1_126 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_7_CLKBUF1_37 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_19_CLKBUF1_2 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_10_DFFPOSX1_30 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_43_DFFSR_29 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_32_DFFSR_69 BUFX2_98/A DFFSR_32/S FILL
XFILL_6_CLKBUF1_40 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_49_DFFSR_125 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_5_CLKBUF1_43 AND2X2_38/B DFFSR_23/S FILL
XNAND3X1_162 AOI21X1_10/B AOI21X1_10/A AOI21X1_10/C BUFX2_8/gnd AOI21X1_20/B DFFSR_51/S
+ NAND3X1
XCLKBUF1_40 BUFX2_6/Y OR2X2_6/gnd CLKBUF1_40/Y DFFSR_92/S CLKBUF1
XFILL_39_DFFSR_128 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_16_DFFSR_19 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_2_DFFSR_204 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_4_CLKBUF1_46 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_3_BUFX2_54 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_29_DFFSR_131 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_43_DFFSR_235 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_3_CLKBUF1_49 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_19_DFFSR_134 INVX1_1/gnd DFFSR_53/S FILL
XFILL_20_DFFPOSX1_19 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_33_DFFSR_238 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_6_0_2 BUFX2_7/gnd DFFSR_216/S FILL
XNOR2X1_16 NOR2X1_16/A OAI21X1_4/Y BUFX2_79/A NOR2X1_16/Y DFFSR_7/S NOR2X1
XFILL_48_DFFSR_3 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_23_DFFSR_241 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_4_NAND3X1_222 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_51_DFFSR_36 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_4_XNOR2X1_4 BUFX2_98/A DFFSR_6/S FILL
XFILL_40_DFFSR_76 BUFX2_79/A DFFSR_7/S FILL
XFILL_4_NOR2X1_13 BUFX2_99/A DFFSR_92/S FILL
XFILL_0_DFFPOSX1_41 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_13_DFFSR_244 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_50_3 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_7_DFFSR_33 BUFX2_98/A DFFSR_32/S FILL
XFILL_24_DFFSR_26 BUFX2_79/A DFFSR_6/S FILL
XFILL_13_DFFSR_66 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_5_DFFSR_131 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_46_DFFSR_162 BUFX2_99/A DFFSR_92/S FILL
XFILL_5_NAND3X1_156 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_9_DFFSR_238 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_53_2_0 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_16_XOR2X1_13 INVX1_1/gnd DFFSR_97/S FILL
XFILL_36_DFFSR_165 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_3_INVX1_5 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_50_DFFSR_269 INVX1_67/gnd DFFSR_201/S FILL
XFILL_0_XOR2X1_3 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_26_DFFSR_168 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_2_INVX1_215 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_40_DFFSR_272 INVX1_3/gnd DFFSR_23/S FILL
XFILL_51_4_1 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_48_DFFSR_83 INVX1_3/gnd DFFSR_79/S FILL
XFILL_16_DFFSR_171 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_30_DFFSR_275 BUFX2_99/A DFFSR_92/S FILL
XFILL_8_AOI22X1_3 INVX1_1/gnd DFFSR_97/S FILL
XFILL_4_INVX1_27 BUFX2_99/A DFFSR_7/S FILL
XFILL_20_DFFSR_278 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_49_6_2 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_4_DFFSR_80 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_32_DFFSR_33 BUFX2_98/A DFFSR_32/S FILL
XFILL_19_DFFPOSX1_49 BUFX2_99/A DFFSR_92/S FILL
XFILL_21_DFFSR_73 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_2_XOR2X1_10 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_1_NOR2X1_50 INVX1_39/gnd DFFSR_34/S FILL
XNAND3X1_126 DFFSR_208/D BUFX2_28/Y NOR2X1_31/Y DFFSR_62/gnd NAND3X1_126/Y DFFSR_62/S
+ NAND3X1
XFILL_4_CLKBUF1_10 INVX1_67/gnd DFFSR_201/S FILL
XFILL_2_DFFSR_168 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_3_BUFX2_18 BUFX2_98/A DFFSR_32/S FILL
XFILL_3_CLKBUF1_13 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_43_DFFSR_199 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_6_DFFSR_275 BUFX2_99/A DFFSR_92/S FILL
XFILL_6_OAI21X1_108 INVX1_1/gnd DFFSR_53/S FILL
XFILL_2_CLKBUF1_16 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_33_DFFSR_202 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_14_DFFSR_1 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_23_DFFSR_205 INVX1_3/gnd DFFSR_79/S FILL
XFILL_4_NAND3X1_186 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_1_CLKBUF1_19 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_40_DFFSR_40 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_1_INVX1_74 BUFX2_99/A DFFSR_92/S FILL
XFILL_29_DFFSR_80 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_17_5_0 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_0_CLKBUF1_22 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_13_DFFSR_208 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_16_CLKBUF1_3 BUFX2_98/A DFFSR_6/S FILL
XFILL_13_DFFSR_30 BUFX2_98/A DFFSR_32/S FILL
XFILL_0_BUFX2_65 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_46_DFFSR_126 BUFX2_99/A DFFSR_7/S FILL
XFILL_5_NAND3X1_120 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_9_DFFSR_202 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_36_DFFSR_129 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_50_DFFSR_233 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_26_DFFSR_132 INVX1_3/gnd DFFSR_79/S FILL
XFILL_2_INVX1_179 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_40_DFFSR_236 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_37_DFFSR_87 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_48_DFFSR_47 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_16_DFFSR_135 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_30_DFFSR_239 INVX1_39/gnd DFFSR_54/S FILL
XFILL_20_DFFSR_242 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_21_DFFSR_37 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_4_DFFSR_44 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_10_DFFSR_77 BUFX2_98/A DFFSR_32/S FILL
XFILL_19_DFFPOSX1_13 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_1_NOR2X1_14 INVX1_1/gnd DFFSR_97/S FILL
XFILL_10_DFFSR_245 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_3_NAND3X1_216 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_2_DFFSR_132 INVX1_3/gnd DFFSR_79/S FILL
XFILL_27_DFFPOSX1_1 INVX1_39/gnd DFFSR_34/S FILL
XFILL_55_8 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_14_XOR2X1_7 BUFX2_98/A DFFSR_6/S FILL
XFILL_43_DFFSR_163 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_45_DFFSR_94 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_13_XOR2X1_14 INVX1_1/gnd DFFSR_53/S FILL
XFILL_6_DFFSR_239 INVX1_39/gnd DFFSR_54/S FILL
XFILL_26_DFFPOSX1_4 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_33_DFFSR_166 AND2X2_38/B DFFSR_59/S FILL
XFILL_27_0_0 INVX1_3/gnd DFFSR_79/S FILL
XFILL_47_DFFSR_270 INVX1_39/gnd DFFSR_54/S FILL
XFILL_25_DFFPOSX1_7 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_23_DFFSR_169 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_6_AND2X2_3 INVX1_1/gnd DFFSR_53/S FILL
XFILL_4_NAND3X1_150 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_1_DFFSR_91 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_1_INVX1_38 AND2X2_38/B DFFSR_23/S FILL
XFILL_37_DFFSR_273 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_29_DFFSR_44 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_18_DFFSR_84 BUFX2_99/A DFFSR_7/S FILL
XFILL_13_DFFSR_172 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_27_DFFSR_276 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_5_AOI22X1_4 BUFX2_99/A DFFSR_92/S FILL
XOAI21X1_108 DFFSR_91/S INVX1_206/Y NAND2X1_139/Y INVX1_1/gnd DFFSR_280/D DFFSR_53/S
+ OAI21X1
XFILL_25_2_1 AND2X2_38/B DFFSR_23/S FILL
XFILL_9_DFFPOSX1_24 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_7_1_0 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_17_DFFSR_279 BUFX2_99/A DFFSR_7/S FILL
XFILL_0_BUFX2_29 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_23_4_2 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_9_DFFSR_166 AND2X2_38/B DFFSR_59/S FILL
XFILL_5_3_1 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_18_DFFPOSX1_43 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_50_DFFSR_197 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_2_INVX1_143 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_40_DFFSR_200 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_5_AND2X2_10 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_9_DFFSR_98 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_26_DFFSR_91 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_37_DFFSR_51 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_48_DFFSR_11 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_2_NAND3X1_246 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_3_DFFSR_276 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_3_5_2 INVX1_67/gnd DFFSR_175/S FILL
XFILL_30_DFFSR_203 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_20_DFFSR_206 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_10_DFFSR_41 BUFX2_98/A DFFSR_6/S FILL
XFILL_5_OAI21X1_102 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_10_DFFSR_209 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_3_NAND3X1_180 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_13_CLKBUF1_4 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_43_DFFSR_127 BUFX2_99/A DFFSR_92/S FILL
XFILL_45_DFFSR_58 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_34_DFFSR_98 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_6_DFFSR_203 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_33_DFFSR_130 BUFX2_79/A DFFSR_6/S FILL
XFILL_47_DFFSR_234 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_23_DFFSR_133 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_4_NAND3X1_114 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_1_DFFSR_55 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_37_DFFSR_237 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_18_DFFSR_48 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_13_DFFSR_136 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_5_BUFX2_83 BUFX2_79/A DFFSR_7/S FILL
XFILL_15_5 INVX1_39/gnd DFFSR_54/S FILL
XFILL_27_DFFSR_240 INVX1_39/gnd DFFSR_34/S FILL
XFILL_8_XNOR2X1_3 INVX1_1/gnd DFFSR_97/S FILL
XFILL_6_NAND2X1_150 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_17_DFFSR_243 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_26_DFFSR_4 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_9_DFFSR_130 BUFX2_79/A DFFSR_6/S FILL
XFILL_50_DFFSR_161 INVX1_67/gnd DFFSR_175/S FILL
XFILL_40_DFFSR_164 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_2_INVX1_107 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_37_DFFSR_15 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_26_DFFSR_55 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_9_DFFSR_62 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_15_DFFSR_95 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_2_NAND3X1_210 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_10_XOR2X1_15 BUFX2_99/A DFFSR_7/S FILL
XFILL_3_DFFSR_240 INVX1_39/gnd DFFSR_34/S FILL
XFILL_30_DFFSR_167 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_44_DFFSR_271 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_20_DFFSR_170 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_34_DFFSR_274 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_10_DFFSR_173 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_24_DFFSR_277 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_2_AOI22X1_5 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_15_DFFPOSX1_1 INVX1_39/gnd DFFSR_34/S FILL
XFILL_3_NAND3X1_144 AND2X2_38/B DFFSR_59/S FILL
XFILL_5_NOR2X1_49 AND2X2_38/B DFFSR_59/S FILL
XFILL_14_DFFSR_280 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_14_DFFPOSX1_4 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_13_DFFPOSX1_7 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_8_DFFPOSX1_18 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_45_DFFSR_22 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_5_NAND2X1_180 INVX1_1/gnd DFFSR_97/S FILL
XFILL_6_DFFSR_167 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_34_DFFSR_62 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_47_DFFSR_198 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_37_DFFSR_201 INVX1_67/gnd DFFSR_201/S FILL
XFILL_1_DFFSR_19 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_18_DFFSR_12 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_2_AND2X2_11 BUFX2_99/A DFFSR_7/S FILL
XBUFX2_87 BUFX2_87/A INVX1_1/gnd BUFX2_87/Y DFFSR_53/S BUFX2
XFILL_13_DFFSR_100 INVX1_1/gnd DFFSR_97/S FILL
XFILL_0_DFFSR_277 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_5_BUFX2_47 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_17_DFFPOSX1_37 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_27_DFFSR_204 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_6_NAND2X1_114 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_2_INVX1_2 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_17_DFFSR_207 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_1_NAND3X1_240 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_20_CLKBUF1_2 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_42_DFFSR_69 BUFX2_98/A DFFSR_32/S FILL
XNAND2X1_150 NAND2X1_149/B INVX1_208/Y DFFSR_1/gnd AOI21X1_51/A DFFSR_1/S NAND2X1
XFILL_50_DFFSR_125 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_10_CLKBUF1_5 BUFX2_99/A DFFSR_92/S FILL
XFILL_27_DFFPOSX1_26 AND2X2_38/B DFFSR_23/S FILL
XFILL_8_AOI21X1_42 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_40_DFFSR_128 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_7_AOI21X1_45 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_26_DFFSR_19 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_9_DFFSR_26 BUFX2_79/A DFFSR_6/S FILL
XFILL_15_DFFSR_59 AND2X2_38/B DFFSR_59/S FILL
XFILL_2_NAND3X1_174 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_3_DFFSR_204 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_30_DFFSR_131 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_24_5_0 AND2X2_38/B DFFSR_59/S FILL
XFILL_2_BUFX2_94 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_6_AOI21X1_48 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_44_DFFSR_235 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_20_DFFSR_134 INVX1_1/gnd DFFSR_53/S FILL
XFILL_7_DFFPOSX1_48 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_34_DFFSR_238 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_5_AOI21X1_51 DFFSR_1/gnd DFFSR_81/S FILL
XAOI21X1_48 AOI21X1_48/A AOI21X1_48/B BUFX2_39/Y DFFSR_62/gnd AOI21X1_48/Y DFFSR_62/S
+ AOI21X1
XFILL_10_DFFSR_137 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_4_AOI21X1_54 AND2X2_38/B DFFSR_59/S FILL
XFILL_24_DFFSR_241 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_5_XNOR2X1_4 BUFX2_98/A DFFSR_6/S FILL
XFILL_50_DFFSR_76 BUFX2_79/A DFFSR_7/S FILL
XFILL_5_NOR2X1_13 BUFX2_99/A DFFSR_92/S FILL
XFILL_3_NAND3X1_108 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_3_AOI21X1_57 INVX1_67/gnd DFFSR_201/S FILL
XFILL_4_6_0 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_14_DFFSR_244 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_37_5 BUFX2_99/A DFFSR_92/S FILL
XFILL_2_AOI21X1_60 BUFX2_79/A DFFSR_7/S FILL
XFILL_6_DFFSR_73 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_5_NAND2X1_144 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_23_DFFSR_66 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_34_DFFSR_26 BUFX2_79/A DFFSR_6/S FILL
XFILL_6_DFFSR_131 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_1_AOI21X1_63 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_47_DFFSR_162 BUFX2_99/A DFFSR_92/S FILL
XFILL_0_AOI21X1_66 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_37_DFFSR_165 BUFX2_72/gnd DFFSR_201/S FILL
XBUFX2_51 INVX1_59/Y OR2X2_3/gnd DFFSR_5/R DFFSR_4/S BUFX2
XFILL_0_DFFSR_241 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_5_BUFX2_11 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_27_DFFSR_168 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_41_DFFSR_272 INVX1_3/gnd DFFSR_23/S FILL
XFILL_3_INVX1_215 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_17_DFFSR_171 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_8_OAI21X1_90 BUFX2_98/A DFFSR_32/S FILL
XFILL_31_DFFSR_275 BUFX2_99/A DFFSR_92/S FILL
XFILL_9_AOI22X1_3 INVX1_1/gnd DFFSR_97/S FILL
XFILL_1_NAND3X1_204 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_7_OAI21X1_93 OR2X2_2/gnd DFFSR_175/S FILL
XOAI21X1_1 INVX1_9/Y OAI21X1_4/B OAI21X1_1/C BUFX2_79/A NOR2X1_6/B DFFSR_7/S OAI21X1
XFILL_21_DFFSR_278 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_3_INVX1_67 INVX1_67/gnd DFFSR_201/S FILL
XFILL_42_DFFSR_33 BUFX2_98/A DFFSR_32/S FILL
XFILL_31_DFFSR_73 OR2X2_1/gnd DFFSR_51/S FILL
XNAND2X1_114 INVX1_180/Y AND2X2_40/A OR2X2_4/gnd NAND2X1_114/Y DFFSR_32/S NAND2X1
XFILL_3_XOR2X1_10 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_2_NOR2X1_50 INVX1_39/gnd DFFSR_34/S FILL
XFILL_6_OAI21X1_96 AND2X2_38/B DFFSR_59/S FILL
XFILL_34_0_0 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_5_OAI21X1_99 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_15_DFFSR_23 AND2X2_38/B DFFSR_23/S FILL
XOAI21X1_96 BUFX2_55/Y INVX1_193/Y OAI21X1_96/C AND2X2_38/B DFFSR_268/D DFFSR_59/S
+ OAI21X1
XFILL_2_NAND3X1_138 INVX1_67/gnd DFFSR_201/S FILL
XFILL_3_DFFSR_168 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_2_BUFX2_58 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_6_AOI21X1_12 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_44_DFFSR_199 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_32_2_1 INVX1_1/gnd DFFSR_97/S FILL
XFILL_7_DFFPOSX1_12 AND2X2_38/B DFFSR_23/S FILL
XFILL_7_DFFSR_275 BUFX2_99/A DFFSR_92/S FILL
XFILL_5_AOI21X1_15 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_4_NAND2X1_174 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_6_NOR3X1_4 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_34_DFFSR_202 NOR3X1_6/gnd DFFSR_91/S FILL
XAOI21X1_12 AOI21X1_12/A AOI21X1_12/B AOI21X1_12/C DFFSR_1/gnd OAI21X1_40/B DFFSR_1/S
+ AOI21X1
XFILL_10_DFFSR_101 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_38_DFFSR_7 BUFX2_79/A DFFSR_7/S FILL
XFILL_3_DFFPOSX1_1 INVX1_39/gnd DFFSR_34/S FILL
XFILL_4_AOI21X1_18 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_24_DFFSR_205 INVX1_3/gnd DFFSR_79/S FILL
XFILL_50_DFFSR_40 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_30_4_2 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_39_DFFSR_80 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_3_AOI21X1_21 INVX1_39/gnd DFFSR_54/S FILL
XFILL_2_DFFPOSX1_4 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_14_DFFSR_208 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_1_DFFPOSX1_7 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_16_DFFPOSX1_31 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_2_AOI21X1_24 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_17_CLKBUF1_3 BUFX2_98/A DFFSR_6/S FILL
XFILL_6_DFFSR_37 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_5_NAND2X1_108 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_12_DFFSR_70 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_23_DFFSR_30 BUFX2_98/A DFFSR_32/S FILL
XFILL_1_AOI21X1_27 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_0_NAND3X1_234 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_47_DFFSR_126 BUFX2_99/A DFFSR_7/S FILL
XFILL_0_AOI21X1_30 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_37_DFFSR_129 XOR2X1_1/gnd DFFSR_151/S FILL
XBUFX2_15 NOR2X1_7/Y DFFSR_8/gnd BUFX2_15/Y DFFSR_8/S BUFX2
XFILL_0_DFFSR_205 INVX1_3/gnd DFFSR_79/S FILL
XFILL_27_DFFSR_132 INVX1_3/gnd DFFSR_79/S FILL
XFILL_3_INVX1_179 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_26_DFFPOSX1_20 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_41_DFFSR_236 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_47_DFFSR_87 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_17_DFFSR_135 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_31_DFFSR_239 INVX1_39/gnd DFFSR_54/S FILL
XFILL_8_OAI21X1_54 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_1_NAND3X1_168 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_6_NAND2X1_75 INVX1_3/gnd DFFSR_79/S FILL
XFILL_7_OAI21X1_57 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_21_DFFSR_242 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_31_DFFSR_37 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_3_DFFSR_84 BUFX2_99/A DFFSR_7/S FILL
XFILL_3_INVX1_31 INVX1_1/gnd DFFSR_53/S FILL
XFILL_20_DFFSR_77 BUFX2_98/A DFFSR_32/S FILL
XFILL_2_NOR2X1_14 INVX1_1/gnd DFFSR_97/S FILL
XFILL_6_DFFPOSX1_42 INVX1_39/gnd DFFSR_34/S FILL
XFILL_5_NAND2X1_78 AND2X2_38/B DFFSR_23/S FILL
XFILL_6_OAI21X1_60 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_11_DFFSR_245 DFFSR_34/gnd DFFSR_34/S FILL
XNAND2X1_75 INVX1_135/A AND2X2_34/B INVX1_3/gnd NAND2X1_77/A DFFSR_79/S NAND2X1
XFILL_5_OAI21X1_63 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_4_NAND2X1_81 DFFSR_34/gnd DFFSR_34/S FILL
XOAI21X1_60 OAI21X1_36/C XOR2X1_4/A AOI22X1_23/A OR2X2_1/gnd XNOR2X1_1/A DFFSR_51/S
+ OAI21X1
XFILL_2_NAND3X1_102 INVX1_3/gnd DFFSR_23/S FILL
XFILL_4_OAI21X1_66 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_3_NAND2X1_84 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_3_DFFSR_132 INVX1_3/gnd DFFSR_79/S FILL
XFILL_2_BUFX2_22 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_44_DFFSR_163 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_2_NAND2X1_87 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_3_OAI21X1_69 INVX1_3/gnd DFFSR_23/S FILL
XFILL_14_XOR2X1_14 INVX1_1/gnd DFFSR_53/S FILL
XFILL_7_DFFSR_239 INVX1_39/gnd DFFSR_54/S FILL
XFILL_4_NAND2X1_138 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_34_DFFSR_166 AND2X2_38/B DFFSR_59/S FILL
XFILL_12_NOR3X1_1 INVX1_3/gnd DFFSR_79/S FILL
XFILL_2_OAI21X1_72 INVX1_3/gnd DFFSR_23/S FILL
XFILL_1_NAND2X1_90 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_48_DFFSR_270 INVX1_39/gnd DFFSR_54/S FILL
XFILL_24_DFFSR_169 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_0_NAND2X1_93 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_1_OAI21X1_75 INVX1_39/gnd DFFSR_54/S FILL
XFILL_38_DFFSR_273 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_39_DFFSR_44 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_28_DFFSR_84 BUFX2_99/A DFFSR_7/S FILL
XFILL_0_INVX1_216 INVX1_1/gnd DFFSR_97/S FILL
XFILL_0_INVX1_78 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_14_DFFSR_172 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_0_OAI21X1_78 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_28_DFFSR_276 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_6_AOI22X1_4 BUFX2_99/A DFFSR_92/S FILL
XFILL_18_DFFSR_279 BUFX2_99/A DFFSR_7/S FILL
XFILL_25_DFFPOSX1_50 INVX1_1/gnd DFFSR_53/S FILL
XFILL_12_DFFSR_34 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_0_XOR2X1_11 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_0_NAND3X1_198 DFFSR_62/gnd DFFSR_62/S FILL
XDFFSR_279 BUFX2_77/A DFFSR_2/CLK DFFSR_274/R DFFSR_7/S DFFSR_279/D BUFX2_99/A DFFSR_7/S
+ DFFSR
XFILL_0_DFFSR_169 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_25_DFFSR_1 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_9_OAI21X1_15 INVX1_3/gnd DFFSR_79/S FILL
XFILL_3_INVX1_143 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_41_DFFSR_200 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_6_AND2X2_10 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_36_DFFSR_91 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_47_DFFSR_51 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_4_DFFSR_276 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_8_OAI21X1_18 INVX1_39/gnd DFFSR_34/S FILL
XFILL_31_DFFSR_203 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_1_NAND3X1_132 AND2X2_38/B DFFSR_23/S FILL
XFILL_6_NAND2X1_39 BUFX2_98/A DFFSR_6/S FILL
XFILL_7_OAI21X1_21 AND2X2_38/B DFFSR_59/S FILL
XFILL_21_DFFSR_206 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_3_DFFSR_48 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_20_DFFSR_41 BUFX2_98/A DFFSR_6/S FILL
XFILL_6_OAI21X1_24 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_5_NAND2X1_42 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_11_DFFSR_209 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_3_NAND2X1_168 BUFX2_79/A DFFSR_6/S FILL
XNAND2X1_39 DFFSR_242/D NOR2X1_34/Y BUFX2_98/A OAI21X1_10/C DFFSR_6/S NAND2X1
XFILL_4_NAND2X1_45 INVX1_39/gnd DFFSR_34/S FILL
XFILL_5_OAI21X1_27 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_14_CLKBUF1_4 OR2X2_3/gnd DFFSR_60/S FILL
XOAI21X1_24 INVX1_139/A NOR2X1_65/Y INVX1_138/A DFFSR_34/gnd NAND2X1_64/B DFFSR_1/S
+ OAI21X1
XFILL_3_NAND2X1_48 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_4_OAI21X1_30 DFFSR_1/gnd DFFSR_81/S FILL
XDFFPOSX1_42 AND2X2_35/B CLKBUF1_47/Y NOR3X1_6/Y INVX1_39/gnd DFFSR_34/S DFFPOSX1
XFILL_44_DFFSR_127 BUFX2_99/A DFFSR_92/S FILL
XFILL_15_DFFPOSX1_25 BUFX2_79/A DFFSR_6/S FILL
XFILL_2_NAND2X1_51 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_3_OAI21X1_33 INVX1_3/gnd DFFSR_79/S FILL
XFILL_44_DFFSR_98 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_7_DFFSR_203 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_34_DFFSR_130 BUFX2_79/A DFFSR_6/S FILL
XFILL_4_NAND2X1_102 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_1_NAND2X1_54 AND2X2_38/B DFFSR_59/S FILL
XFILL_2_OAI21X1_36 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_48_DFFSR_234 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_24_DFFSR_133 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_5_AND2X2_7 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_0_NAND2X1_57 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_38_DFFSR_237 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_1_OAI21X1_39 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_28_DFFSR_48 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_17_DFFSR_88 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_0_DFFSR_95 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_0_INVX1_42 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_0_INVX1_180 BUFX2_98/A DFFSR_6/S FILL
XFILL_0_CLKBUF1_1 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_14_DFFSR_136 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_19_2 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_0_OAI21X1_42 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_28_DFFSR_240 INVX1_39/gnd DFFSR_34/S FILL
XFILL_9_XNOR2X1_3 INVX1_1/gnd DFFSR_97/S FILL
XFILL_18_DFFSR_243 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_25_DFFPOSX1_14 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_0_NAND3X1_162 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_8_AOI22X1_11 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_31_5_0 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_9_NAND3X1_217 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_7_AOI22X1_14 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_51_DFFSR_161 INVX1_67/gnd DFFSR_175/S FILL
XFILL_5_DFFPOSX1_36 OR2X2_2/gnd DFFSR_175/S FILL
XDFFSR_243 INVX1_82/A CLKBUF1_11/Y BUFX2_67/Y DFFSR_151/S DFFSR_235/Q BUFX2_7/gnd
+ DFFSR_151/S DFFSR
XFILL_0_DFFSR_133 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_6_AOI22X1_17 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_41_DFFSR_164 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_3_INVX1_107 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_47_DFFSR_15 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_36_DFFSR_55 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_25_DFFSR_95 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_11_XOR2X1_15 BUFX2_99/A DFFSR_7/S FILL
XFILL_5_AOI22X1_20 INVX1_39/gnd DFFSR_34/S FILL
XFILL_4_DFFSR_240 INVX1_39/gnd DFFSR_34/S FILL
XFILL_31_DFFSR_167 OR2X2_2/gnd DFFSR_216/S FILL
XAOI22X1_17 BUFX2_56/Y INVX1_145/A AND2X2_35/A INVX1_135/A NOR3X1_6/gnd INVX1_139/A
+ DFFSR_79/S AOI22X1
XFILL_45_DFFSR_271 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_4_AOI22X1_23 INVX1_39/gnd DFFSR_34/S FILL
XFILL_21_DFFSR_170 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_35_DFFSR_274 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_3_DFFSR_12 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_3_AOI22X1_26 INVX1_1/gnd DFFSR_97/S FILL
XFILL_3_NAND2X1_132 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_11_DFFSR_173 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_25_DFFSR_277 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_3_AOI22X1_5 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_2_AOI22X1_29 INVX1_1/gnd DFFSR_53/S FILL
XFILL_6_NOR2X1_49 AND2X2_38/B DFFSR_59/S FILL
XFILL_15_DFFSR_280 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_3_NAND2X1_12 INVX1_3/gnd DFFSR_79/S FILL
XFILL_2_NAND2X1_15 BUFX2_99/A DFFSR_92/S FILL
XFILL_1_OAI21X1_114 AND2X2_38/B DFFSR_59/S FILL
XFILL_44_DFFSR_62 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_7_DFFSR_167 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_24_DFFPOSX1_44 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_1_NAND2X1_18 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_48_DFFSR_198 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_8_NAND3X1_74 INVX1_1/gnd DFFSR_97/S FILL
XFILL_38_DFFSR_201 INVX1_67/gnd DFFSR_201/S FILL
XFILL_0_NAND2X1_21 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_8_NAND3X1_247 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_28_DFFSR_12 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_17_DFFSR_52 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_0_DFFSR_59 AND2X2_38/B DFFSR_59/S FILL
XFILL_0_INVX1_144 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_3_AND2X2_11 BUFX2_99/A DFFSR_7/S FILL
XFILL_1_DFFSR_277 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_7_NAND3X1_77 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_4_BUFX2_87 INVX1_1/gnd DFFSR_53/S FILL
XFILL_14_DFFSR_100 INVX1_1/gnd DFFSR_97/S FILL
XFILL_28_DFFSR_204 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_6_NAND3X1_80 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_41_0_0 BUFX2_98/A DFFSR_32/S FILL
XFILL_18_DFFSR_207 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_5_NAND3X1_83 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_0_NAND3X1_126 DFFSR_62/gnd DFFSR_62/S FILL
XNAND3X1_80 NOR2X1_38/Y NOR2X1_39/Y NOR2X1_40/Y NOR3X1_6/gnd XOR2X1_9/B DFFSR_91/S
+ NAND3X1
XFILL_16_DFFSR_8 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_4_NAND3X1_86 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_39_2_1 BUFX2_79/A DFFSR_6/S FILL
XFILL_11_CLKBUF1_5 BUFX2_99/A DFFSR_92/S FILL
XFILL_3_NAND3X1_89 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_2_NAND2X1_162 BUFX2_72/gnd DFFSR_201/S FILL
XDFFSR_207 DFFSR_207/Q CLKBUF1_20/Y BUFX2_66/Y DFFSR_62/S DFFSR_199/Q DFFSR_62/gnd
+ DFFSR_62/S DFFSR
XFILL_41_DFFSR_128 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_2_NAND3X1_92 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_36_DFFSR_19 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_8_DFFSR_66 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_14_DFFSR_99 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_25_DFFSR_59 AND2X2_38/B DFFSR_59/S FILL
XFILL_4_DFFSR_204 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_37_4_2 BUFX2_99/A DFFSR_7/S FILL
XFILL_31_DFFSR_131 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_1_NAND3X1_95 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_45_DFFSR_235 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_0_BUFX2_9 AND2X2_38/B DFFSR_59/S FILL
XFILL_21_DFFSR_134 INVX1_1/gnd DFFSR_53/S FILL
XFILL_0_NAND3X1_98 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_35_DFFSR_238 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_14_DFFPOSX1_19 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_11_DFFSR_137 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_25_DFFSR_241 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_6_XNOR2X1_4 BUFX2_98/A DFFSR_6/S FILL
XFILL_6_NOR2X1_13 BUFX2_99/A DFFSR_92/S FILL
XFILL_24_7 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_37_DFFSR_4 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_15_DFFSR_244 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_10_OAI22X1_17 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_33_DFFSR_66 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_44_DFFSR_26 BUFX2_79/A DFFSR_6/S FILL
XFILL_7_DFFSR_131 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_48_DFFSR_162 BUFX2_99/A DFFSR_92/S FILL
XFILL_9_OAI22X1_20 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_8_NAND3X1_38 BUFX2_98/A DFFSR_32/S FILL
XFILL_38_DFFSR_165 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_8_NAND3X1_211 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_17_DFFSR_16 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_0_INVX1_108 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_0_DFFSR_23 AND2X2_38/B DFFSR_23/S FILL
XFILL_1_DFFSR_241 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_4_BUFX2_51 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_8_OAI22X1_23 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_7_NAND3X1_41 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_28_DFFSR_168 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_4_DFFPOSX1_30 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_42_DFFSR_272 INVX1_3/gnd DFFSR_23/S FILL
XFILL_6_NAND3X1_44 BUFX2_99/A DFFSR_7/S FILL
XFILL_4_INVX1_215 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_7_OAI22X1_26 INVX1_39/gnd DFFSR_54/S FILL
XFILL_18_DFFSR_171 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_5_NAND3X1_47 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_32_DFFSR_275 BUFX2_99/A DFFSR_92/S FILL
XXOR2X1_13 XOR2X1_13/A INVX1_217/A INVX1_1/gnd XOR2X1_13/Y DFFSR_97/S XOR2X1
XFILL_6_OAI22X1_29 INVX1_3/gnd DFFSR_79/S FILL
XNAND3X1_44 NAND2X1_22/Y NAND3X1_41/Y AND2X2_11/Y BUFX2_99/A NOR2X1_23/A DFFSR_7/S
+ NAND3X1
XFILL_0_AOI22X1_6 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_22_DFFSR_278 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_4_NAND3X1_50 BUFX2_98/A DFFSR_6/S FILL
XFILL_41_DFFSR_73 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_5_OAI22X1_32 INVX1_39/gnd DFFSR_54/S FILL
XFILL_4_XOR2X1_10 OR2X2_1/gnd DFFSR_59/S FILL
XOAI22X1_29 INVX1_71/Y OAI22X1_41/B INVX1_72/Y OAI22X1_41/D INVX1_3/gnd NOR2X1_38/A
+ DFFSR_79/S OAI22X1
XFILL_3_NOR2X1_50 INVX1_39/gnd DFFSR_34/S FILL
XFILL_13_DFFPOSX1_49 BUFX2_99/A DFFSR_92/S FILL
XFILL_3_NAND3X1_53 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_4_OAI22X1_35 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_2_NAND2X1_126 OR2X2_2/gnd DFFSR_175/S FILL
XDFFSR_171 DFFSR_187/D CLKBUF1_29/Y BUFX2_61/Y DFFSR_81/S DFFSR_163/Q BUFX2_8/gnd
+ DFFSR_81/S DFFSR
XFILL_2_NAND3X1_56 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_3_OAI22X1_38 AND2X2_38/B DFFSR_23/S FILL
XFILL_8_DFFSR_30 BUFX2_98/A DFFSR_32/S FILL
XFILL_14_DFFSR_63 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_25_DFFSR_23 AND2X2_38/B DFFSR_23/S FILL
XFILL_4_DFFSR_168 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_1_BUFX2_98 BUFX2_79/A DFFSR_7/S FILL
XFILL_1_NAND3X1_59 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_2_OAI22X1_41 INVX1_39/gnd DFFSR_54/S FILL
XFILL_45_DFFSR_199 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_0_NAND3X1_62 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_8_DFFSR_275 BUFX2_99/A DFFSR_92/S FILL
XFILL_1_OAI22X1_44 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_35_DFFSR_202 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_0_OAI21X1_108 INVX1_1/gnd DFFSR_53/S FILL
XFILL_0_AND2X2_12 BUFX2_98/A DFFSR_32/S FILL
XFILL_23_DFFPOSX1_38 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_11_DFFSR_101 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_0_OAI22X1_47 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_25_DFFSR_205 INVX1_3/gnd DFFSR_79/S FILL
XFILL_49_DFFSR_80 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_7_NAND3X1_241 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_15_DFFSR_208 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_18_CLKBUF1_3 BUFX2_98/A DFFSR_6/S FILL
XINVX1_64 INVX1_64/A DFFSR_46/gnd INVX1_64/Y DFFSR_62/S INVX1
XFILL_22_DFFSR_70 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_33_DFFSR_30 BUFX2_98/A DFFSR_32/S FILL
XFILL_5_DFFSR_77 BUFX2_98/A DFFSR_32/S FILL
XFILL_48_DFFSR_126 BUFX2_99/A DFFSR_7/S FILL
XFILL_13_0_1 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_38_DFFSR_129 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_8_NAND3X1_175 NOR3X1_6/gnd DFFSR_91/S FILL
XINVX1_182 DFFSR_2/D BUFX2_77/gnd INVX1_182/Y DFFSR_5/S INVX1
XFILL_4_BUFX2_15 DFFSR_8/gnd DFFSR_8/S FILL
XCLKBUF1_3 BUFX2_6/Y BUFX2_98/A CLKBUF1_3/Y DFFSR_6/S CLKBUF1
XFILL_1_DFFSR_205 INVX1_3/gnd DFFSR_79/S FILL
XFILL_28_DFFSR_132 INVX1_3/gnd DFFSR_79/S FILL
XFILL_9_XOR2X1_7 BUFX2_98/A DFFSR_6/S FILL
XFILL_1_NAND2X1_156 AND2X2_38/B DFFSR_59/S FILL
XFILL_11_2_2 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_42_DFFSR_236 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_4_INVX1_179 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_4_DFFSR_7 BUFX2_79/A DFFSR_7/S FILL
XFILL_18_DFFSR_135 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_5_NAND3X1_11 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_32_DFFSR_239 INVX1_39/gnd DFFSR_54/S FILL
XFILL_22_DFFSR_242 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_41_DFFSR_37 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_4_NAND3X1_14 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_2_INVX1_71 BUFX2_79/A DFFSR_6/S FILL
XFILL_30_DFFSR_77 BUFX2_98/A DFFSR_32/S FILL
XFILL_3_NOR2X1_14 INVX1_1/gnd DFFSR_97/S FILL
XFILL_13_DFFPOSX1_13 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_12_DFFSR_245 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_3_NAND3X1_17 BUFX2_99/A DFFSR_7/S FILL
XDFFSR_135 DFFSR_135/Q CLKBUF1_31/Y BUFX2_68/Y DFFSR_208/S BUFX2_88/A DFFSR_62/gnd
+ DFFSR_208/S DFFSR
XFILL_2_NAND3X1_20 BUFX2_99/A DFFSR_7/S FILL
XFILL_14_DFFSR_27 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_4_DFFSR_132 INVX1_3/gnd DFFSR_79/S FILL
XFILL_1_NAND3X1_23 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_1_BUFX2_62 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_45_DFFSR_163 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_0_NAND3X1_26 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_15_XOR2X1_14 INVX1_1/gnd DFFSR_53/S FILL
XFILL_8_DFFSR_239 INVX1_39/gnd DFFSR_54/S FILL
XFILL_35_DFFSR_166 AND2X2_38/B DFFSR_59/S FILL
XFILL_49_DFFSR_270 INVX1_39/gnd DFFSR_54/S FILL
XFILL_0_OAI22X1_11 BUFX2_99/A DFFSR_92/S FILL
XFILL_25_DFFSR_169 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_39_DFFSR_273 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_49_DFFSR_44 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_38_DFFSR_84 BUFX2_99/A DFFSR_7/S FILL
XFILL_1_INVX1_216 INVX1_1/gnd DFFSR_97/S FILL
XFILL_38_5_0 BUFX2_79/A DFFSR_7/S FILL
XFILL_7_NAND3X1_205 INVX1_1/gnd DFFSR_53/S FILL
XFILL_15_DFFSR_172 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_29_DFFSR_276 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_7_AOI22X1_4 BUFX2_99/A DFFSR_92/S FILL
XFILL_3_DFFPOSX1_24 BUFX2_8/gnd DFFSR_51/S FILL
XINVX1_28 INVX1_28/A DFFSR_28/gnd INVX1_28/Y DFFSR_3/S INVX1
XFILL_19_DFFSR_279 BUFX2_99/A DFFSR_7/S FILL
XDFFSR_81 INVX1_5/A CLKBUF1_8/Y DFFSR_1/R DFFSR_81/S INVX1_6/A DFFSR_1/gnd DFFSR_81/S
+ DFFSR
XFILL_5_DFFSR_41 BUFX2_98/A DFFSR_6/S FILL
XFILL_22_DFFSR_34 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_11_DFFSR_74 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_1_XOR2X1_11 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_0_NOR2X1_51 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_8_NAND3X1_139 BUFX2_8/gnd DFFSR_51/S FILL
XINVX1_146 AND2X2_34/B INVX1_3/gnd INVX1_146/Y DFFSR_79/S INVX1
XFILL_12_DFFPOSX1_43 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_1_DFFSR_169 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_49_DFFSR_7 BUFX2_79/A DFFSR_7/S FILL
XFILL_15_XOR2X1_4 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_1_NAND2X1_120 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_42_DFFSR_200 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_7_AND2X2_10 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_46_DFFSR_91 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_5_DFFSR_276 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_32_DFFSR_203 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_22_DFFSR_206 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_2_INVX1_35 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_2_DFFSR_88 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_30_DFFSR_41 BUFX2_98/A DFFSR_6/S FILL
XFILL_19_DFFSR_81 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_12_DFFSR_209 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_22_DFFPOSX1_32 INVX1_67/gnd DFFSR_201/S FILL
XFILL_15_CLKBUF1_4 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_6_NAND3X1_235 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_1_BUFX2_26 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_4_INVX1_9 BUFX2_99/A DFFSR_7/S FILL
XFILL_45_DFFSR_127 BUFX2_99/A DFFSR_92/S FILL
XFILL_8_DFFSR_203 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_35_DFFSR_130 BUFX2_79/A DFFSR_6/S FILL
XFILL_11_NOR3X1_5 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_48_0_0 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_49_DFFSR_234 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_25_DFFSR_133 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_39_DFFSR_237 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_38_DFFSR_48 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_27_DFFSR_88 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_1_INVX1_180 BUFX2_98/A DFFSR_6/S FILL
XFILL_1_CLKBUF1_1 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_15_DFFSR_136 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_7_NAND3X1_169 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_46_2_1 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_29_DFFSR_240 INVX1_39/gnd DFFSR_34/S FILL
XFILL_19_DFFSR_243 BUFX2_7/gnd DFFSR_151/S FILL
XDFFSR_45 DFFSR_61/D DFFSR_45/CLK DFFSR_35/R DFFSR_60/S DFFSR_45/D DFFSR_8/gnd DFFSR_60/S
+ DFFSR
XFILL_0_NAND2X1_150 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_11_DFFSR_38 BUFX2_98/A DFFSR_6/S FILL
XFILL_0_NOR2X1_15 BUFX2_99/A DFFSR_7/S FILL
XFILL_44_4_2 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_8_NAND3X1_103 AND2X2_38/B DFFSR_23/S FILL
XINVX1_110 INVX1_110/A OR2X2_6/gnd INVX1_110/Y DFFSR_53/S INVX1
XFILL_1_DFFSR_133 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_15_DFFSR_5 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_42_DFFSR_164 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_4_INVX1_107 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_46_DFFSR_55 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_35_DFFSR_95 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_12_XOR2X1_15 BUFX2_99/A DFFSR_7/S FILL
XFILL_5_DFFSR_240 INVX1_39/gnd DFFSR_34/S FILL
XFILL_32_DFFSR_167 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_46_DFFSR_271 BUFX2_8/gnd DFFSR_81/S FILL
XAOI22X1_8 NOR3X1_2/Y DFFSR_112/D DFFSR_96/Q NOR3X1_1/Y DFFSR_28/gnd AOI22X1_8/Y DFFSR_3/S
+ AOI22X1
XFILL_22_DFFSR_170 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_2_DFFSR_52 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_36_DFFSR_274 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_19_DFFSR_45 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_6_BUFX2_80 BUFX2_79/A DFFSR_6/S FILL
XFILL_12_DFFSR_173 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_26_DFFSR_277 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_4_AOI22X1_5 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_12_3_0 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_16_DFFSR_280 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_20_CLKBUF1_35 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_6_NAND3X1_199 INVX1_1/gnd DFFSR_97/S FILL
XFILL_10_5_1 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_19_CLKBUF1_38 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_36_DFFSR_1 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_2_DFFPOSX1_18 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_8_DFFSR_167 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_49_DFFSR_198 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_18_CLKBUF1_41 OR2X2_4/gnd DFFSR_3/S FILL
XAND2X2_14 NOR3X1_3/B NOR3X1_3/A DFFSR_46/gnd BUFX2_23/A DFFSR_54/S AND2X2
XNAND3X1_235 NOR2X1_73/Y NAND3X1_235/B NAND3X1_235/C DFFSR_4/gnd AOI21X1_37/B DFFSR_4/S
+ NAND3X1
XFILL_39_DFFSR_201 INVX1_67/gnd DFFSR_201/S FILL
XFILL_17_CLKBUF1_44 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_38_DFFSR_12 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_27_DFFSR_52 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_1_INVX1_144 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_4_AND2X2_11 BUFX2_99/A DFFSR_7/S FILL
XFILL_16_DFFSR_92 BUFX2_99/A DFFSR_92/S FILL
XFILL_2_DFFSR_277 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_15_DFFSR_100 INVX1_1/gnd DFFSR_97/S FILL
XFILL_7_NAND3X1_133 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_29_DFFSR_204 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_16_CLKBUF1_47 BUFX2_98/A DFFSR_32/S FILL
XFILL_11_DFFPOSX1_37 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_0_NAND2X1_114 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_19_DFFSR_207 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_12_CLKBUF1_5 BUFX2_99/A DFFSR_92/S FILL
XFILL_42_DFFSR_128 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_21_DFFPOSX1_26 AND2X2_38/B DFFSR_23/S FILL
XFILL_46_DFFSR_19 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_24_DFFSR_99 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_35_DFFSR_59 AND2X2_38/B DFFSR_59/S FILL
XFILL_5_DFFSR_204 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_32_DFFSR_131 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_46_DFFSR_235 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_5_NAND3X1_229 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_22_DFFSR_134 INVX1_1/gnd DFFSR_53/S FILL
XFILL_2_DFFSR_16 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_36_DFFSR_238 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_1_DFFPOSX1_48 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_12_DFFSR_137 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_6_BUFX2_44 INVX1_3/gnd DFFSR_79/S FILL
XFILL_26_DFFSR_241 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_7_XNOR2X1_4 BUFX2_98/A DFFSR_6/S FILL
XFILL_20_0_1 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_16_DFFSR_244 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_6_NAND3X1_163 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_43_DFFSR_66 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_8_DFFSR_131 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_18_2_2 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_49_DFFSR_162 BUFX2_99/A DFFSR_92/S FILL
XFILL_0_1_1 BUFX2_72/gnd DFFSR_276/S FILL
XNAND3X1_199 INVX1_135/A AOI22X1_25/B AND2X2_37/Y INVX1_1/gnd OAI21X1_78/C DFFSR_97/S
+ NAND3X1
XFILL_39_DFFSR_165 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_27_DFFSR_16 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_1_INVX1_108 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_16_DFFSR_56 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_2_DFFSR_241 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_3_BUFX2_91 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_29_DFFSR_168 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_16_CLKBUF1_11 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_43_DFFSR_272 INVX1_3/gnd DFFSR_23/S FILL
XFILL_19_DFFSR_171 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_15_CLKBUF1_14 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_33_DFFSR_275 BUFX2_99/A DFFSR_92/S FILL
XNOR2X1_53 NOR2X1_53/A NOR2X1_53/B DFFSR_1/gnd NOR2X1_53/Y DFFSR_81/S NOR2X1
XFILL_14_CLKBUF1_17 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_3_DFFSR_4 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_1_AOI22X1_6 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_23_DFFSR_278 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_5_XOR2X1_10 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_13_CLKBUF1_20 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_4_NOR2X1_50 INVX1_39/gnd DFFSR_34/S FILL
XFILL_12_CLKBUF1_23 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_7_OAI21X1_115 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_7_DFFSR_70 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_24_DFFSR_63 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_11_CLKBUF1_26 INVX1_1/gnd DFFSR_53/S FILL
XFILL_35_DFFSR_23 AND2X2_38/B DFFSR_23/S FILL
XFILL_5_DFFSR_168 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_45_5_0 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_10_CLKBUF1_29 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_46_DFFSR_199 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_5_NAND3X1_193 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_9_DFFSR_275 BUFX2_99/A DFFSR_92/S FILL
XFILL_36_DFFSR_202 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_1_OR2X2_4 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_1_DFFPOSX1_12 AND2X2_38/B DFFSR_23/S FILL
XFILL_1_AND2X2_12 BUFX2_98/A DFFSR_32/S FILL
XFILL_12_DFFSR_101 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_26_DFFSR_205 INVX1_3/gnd DFFSR_79/S FILL
XFILL_9_CLKBUF1_32 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_8_CLKBUF1_35 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_16_DFFSR_208 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_27_DFFSR_8 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_6_NAND3X1_127 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_7_CLKBUF1_38 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_19_CLKBUF1_3 BUFX2_98/A DFFSR_6/S FILL
XFILL_10_DFFPOSX1_31 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_32_DFFSR_70 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_43_DFFSR_30 BUFX2_98/A DFFSR_32/S FILL
XFILL_4_INVX1_64 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_6_CLKBUF1_41 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_49_DFFSR_126 BUFX2_99/A DFFSR_7/S FILL
XFILL_5_CLKBUF1_44 DFFSR_1/gnd DFFSR_81/S FILL
XNAND3X1_163 INVX1_152/A OAI21X1_46/C AOI21X1_20/B DFFSR_1/gnd AOI22X1_20/D DFFSR_1/S
+ NAND3X1
XFILL_39_DFFSR_129 XOR2X1_1/gnd DFFSR_151/S FILL
XCLKBUF1_41 BUFX2_1/Y OR2X2_4/gnd DFFSR_92/CLK DFFSR_3/S CLKBUF1
XFILL_16_DFFSR_20 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_4_CLKBUF1_47 BUFX2_98/A DFFSR_32/S FILL
XFILL_2_DFFSR_205 INVX1_3/gnd DFFSR_79/S FILL
XFILL_3_BUFX2_55 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_29_DFFSR_132 INVX1_3/gnd DFFSR_79/S FILL
XFILL_43_DFFSR_236 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_20_DFFPOSX1_20 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_19_DFFSR_135 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_7_NOR3X1_1 INVX1_3/gnd DFFSR_79/S FILL
XFILL_33_DFFSR_239 INVX1_39/gnd DFFSR_54/S FILL
XNOR2X1_17 NOR2X1_17/A NOR2X1_17/B BUFX2_79/A NOR2X1_17/Y DFFSR_6/S NOR2X1
XFILL_48_DFFSR_4 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_23_DFFSR_242 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_4_NAND3X1_223 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_40_DFFSR_77 BUFX2_98/A DFFSR_32/S FILL
XFILL_4_NOR2X1_14 INVX1_1/gnd DFFSR_97/S FILL
XFILL_13_DFFSR_245 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_0_DFFPOSX1_42 INVX1_39/gnd DFFSR_34/S FILL
XFILL_50_4 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_7_DFFSR_34 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_24_DFFSR_27 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_13_DFFSR_67 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_5_DFFSR_132 INVX1_3/gnd DFFSR_79/S FILL
XFILL_5_NAND3X1_157 INVX1_3/gnd DFFSR_23/S FILL
XFILL_46_DFFSR_163 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_53_2_1 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_16_XOR2X1_14 INVX1_1/gnd DFFSR_53/S FILL
XFILL_9_DFFSR_239 INVX1_39/gnd DFFSR_54/S FILL
XFILL_36_DFFSR_166 AND2X2_38/B DFFSR_59/S FILL
XFILL_3_INVX1_6 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_50_DFFSR_270 INVX1_39/gnd DFFSR_54/S FILL
XFILL_0_XOR2X1_4 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_26_DFFSR_169 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_48_DFFSR_84 BUFX2_99/A DFFSR_7/S FILL
XFILL_2_INVX1_216 INVX1_1/gnd DFFSR_97/S FILL
XFILL_40_DFFSR_273 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_51_4_2 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_16_DFFSR_172 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_30_DFFSR_276 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_8_AOI22X1_4 BUFX2_99/A DFFSR_92/S FILL
XFILL_20_DFFSR_279 BUFX2_99/A DFFSR_7/S FILL
XFILL_4_DFFSR_81 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_32_DFFSR_34 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_21_DFFSR_74 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_19_DFFPOSX1_50 INVX1_1/gnd DFFSR_53/S FILL
XFILL_2_XOR2X1_11 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_1_NOR2X1_51 DFFSR_34/gnd DFFSR_34/S FILL
XNAND3X1_127 NAND3X1_127/A NAND3X1_126/Y AOI22X1_16/Y DFFSR_46/gnd NOR2X1_58/B DFFSR_62/S
+ NAND3X1
XFILL_4_CLKBUF1_11 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_2_DFFSR_169 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_3_BUFX2_19 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_43_DFFSR_200 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_3_CLKBUF1_14 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_8_AND2X2_10 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_6_DFFSR_276 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_6_OAI21X1_109 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_19_3_0 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_14_DFFSR_2 BUFX2_79/A DFFSR_7/S FILL
XFILL_2_CLKBUF1_17 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_33_DFFSR_203 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_23_DFFSR_206 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_4_NAND3X1_187 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_1_CLKBUF1_20 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_40_DFFSR_41 BUFX2_98/A DFFSR_6/S FILL
XFILL_1_INVX1_75 BUFX2_98/A DFFSR_6/S FILL
XFILL_29_DFFSR_81 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_17_5_1 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_13_DFFSR_209 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_0_CLKBUF1_23 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_16_CLKBUF1_4 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_13_DFFSR_31 BUFX2_79/A DFFSR_6/S FILL
XFILL_0_BUFX2_66 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_46_DFFSR_127 BUFX2_99/A DFFSR_92/S FILL
XFILL_5_NAND3X1_121 INVX1_1/gnd DFFSR_97/S FILL
XFILL_9_DFFSR_203 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_36_DFFSR_130 BUFX2_79/A DFFSR_6/S FILL
XFILL_50_DFFSR_234 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_26_DFFSR_133 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_10_1 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_48_DFFSR_48 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_2_INVX1_180 BUFX2_98/A DFFSR_6/S FILL
XFILL_40_DFFSR_237 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_37_DFFSR_88 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_2_CLKBUF1_1 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_16_DFFSR_136 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_30_DFFSR_240 INVX1_39/gnd DFFSR_34/S FILL
XFILL_20_DFFSR_243 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_4_DFFSR_45 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_10_DFFSR_78 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_21_DFFSR_38 BUFX2_98/A DFFSR_6/S FILL
XFILL_19_DFFPOSX1_14 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_1_NOR2X1_15 BUFX2_99/A DFFSR_7/S FILL
XFILL_10_DFFSR_246 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_3_NAND3X1_217 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_2_DFFSR_133 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_27_DFFPOSX1_2 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_43_DFFSR_164 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_14_XOR2X1_8 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_55_9 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_45_DFFSR_95 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_26_DFFPOSX1_5 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_6_DFFSR_240 INVX1_39/gnd DFFSR_34/S FILL
XFILL_13_XOR2X1_15 BUFX2_99/A DFFSR_7/S FILL
XFILL_33_DFFSR_167 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_27_0_1 INVX1_3/gnd DFFSR_79/S FILL
XFILL_47_DFFSR_271 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_25_DFFPOSX1_8 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_23_DFFSR_170 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_6_AND2X2_4 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_4_NAND3X1_151 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_37_DFFSR_274 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_18_DFFSR_85 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_29_DFFSR_45 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_1_DFFSR_92 BUFX2_99/A DFFSR_92/S FILL
XFILL_1_INVX1_39 INVX1_39/gnd DFFSR_34/S FILL
XFILL_13_DFFSR_173 XOR2X1_1/gnd DFFSR_208/S FILL
XOAI21X1_109 BUFX2_9/Y OR2X2_1/A INVX1_209/Y NOR3X1_6/gnd AOI21X1_61/C DFFSR_79/S
+ OAI21X1
XFILL_27_DFFSR_277 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_5_AOI22X1_5 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_25_2_2 AND2X2_38/B DFFSR_23/S FILL
XFILL_9_DFFPOSX1_25 BUFX2_79/A DFFSR_6/S FILL
XFILL_17_DFFSR_280 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_7_1_1 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_0_BUFX2_30 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_9_DFFSR_167 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_5_3_2 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_18_DFFPOSX1_44 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_50_DFFSR_198 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_40_DFFSR_201 INVX1_67/gnd DFFSR_201/S FILL
XFILL_48_DFFSR_12 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_9_DFFSR_99 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_2_INVX1_144 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_37_DFFSR_52 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_5_AND2X2_11 BUFX2_99/A DFFSR_7/S FILL
XFILL_26_DFFSR_92 BUFX2_99/A DFFSR_92/S FILL
XFILL_3_DFFSR_277 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_16_DFFSR_100 INVX1_1/gnd DFFSR_97/S FILL
XFILL_2_NAND3X1_247 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_30_DFFSR_204 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_20_DFFSR_207 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_10_DFFSR_42 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_5_OAI21X1_103 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_10_DFFSR_210 BUFX2_98/A DFFSR_6/S FILL
XFILL_52_5_0 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_3_NAND3X1_181 INVX1_39/gnd DFFSR_54/S FILL
XFILL_13_CLKBUF1_5 BUFX2_99/A DFFSR_92/S FILL
XFILL_2_DFFSR_1 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_43_DFFSR_128 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_34_DFFSR_99 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_45_DFFSR_59 AND2X2_38/B DFFSR_59/S FILL
XFILL_6_DFFSR_204 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_33_DFFSR_131 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_47_DFFSR_235 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_4_NAND3X1_115 BUFX2_79/A DFFSR_7/S FILL
XFILL_23_DFFSR_134 INVX1_1/gnd DFFSR_53/S FILL
XFILL_37_DFFSR_238 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_1_DFFSR_56 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_18_DFFSR_49 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_13_DFFSR_137 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_5_BUFX2_84 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_27_DFFSR_241 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_8_XNOR2X1_4 BUFX2_98/A DFFSR_6/S FILL
XFILL_32_1 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_0_OR2X2_1 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_6_NAND2X1_151 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_17_DFFSR_244 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_26_DFFSR_5 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_9_DFFSR_131 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_50_DFFSR_162 BUFX2_99/A DFFSR_92/S FILL
XFILL_40_DFFSR_165 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_37_DFFSR_16 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_9_DFFSR_63 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_2_INVX1_108 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_26_DFFSR_56 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_15_DFFSR_96 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_3_DFFSR_241 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_2_NAND3X1_211 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_30_DFFSR_168 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_44_DFFSR_272 INVX1_3/gnd DFFSR_23/S FILL
XFILL_20_DFFSR_171 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_34_DFFSR_275 BUFX2_99/A DFFSR_92/S FILL
XFILL_10_DFFSR_174 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_2_AOI22X1_6 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_24_DFFSR_278 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_15_DFFPOSX1_2 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_6_XOR2X1_10 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_3_NAND3X1_145 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_5_NOR2X1_50 INVX1_39/gnd DFFSR_34/S FILL
XFILL_14_DFFPOSX1_5 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_47_DFFSR_1 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_8_DFFPOSX1_19 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_13_DFFPOSX1_8 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_34_DFFSR_63 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_5_NAND2X1_181 BUFX2_99/A DFFSR_92/S FILL
XFILL_45_DFFSR_23 AND2X2_38/B DFFSR_23/S FILL
XFILL_6_DFFSR_168 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_47_DFFSR_199 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_1_DFFSR_20 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_18_DFFSR_13 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_37_DFFSR_202 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_2_AND2X2_12 BUFX2_98/A DFFSR_32/S FILL
XFILL_13_DFFSR_101 OR2X2_3/gnd DFFSR_4/S FILL
XBUFX2_88 BUFX2_88/A INVX1_3/gnd BUFX2_88/Y DFFSR_23/S BUFX2
XFILL_0_DFFSR_278 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_5_BUFX2_48 AND2X2_38/B DFFSR_59/S FILL
XFILL_17_DFFPOSX1_38 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_27_DFFSR_205 INVX1_3/gnd DFFSR_79/S FILL
XFILL_6_NAND2X1_115 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_2_INVX1_3 INVX1_3/gnd DFFSR_79/S FILL
XFILL_17_DFFSR_208 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_1_NAND3X1_241 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_0_NOR2X1_1 BUFX2_99/A DFFSR_92/S FILL
XFILL_20_CLKBUF1_3 BUFX2_98/A DFFSR_6/S FILL
XFILL_42_DFFSR_70 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_9_AOI21X1_40 INVX1_39/gnd DFFSR_54/S FILL
XNAND2X1_151 DFFSR_81/S NAND2X1_151/B DFFSR_1/gnd AOI21X1_51/B DFFSR_81/S NAND2X1
XFILL_10_CLKBUF1_6 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_50_DFFSR_126 BUFX2_99/A DFFSR_7/S FILL
XFILL_26_3_0 INVX1_3/gnd DFFSR_23/S FILL
XFILL_8_AOI21X1_43 INVX1_3/gnd DFFSR_79/S FILL
XFILL_27_DFFPOSX1_27 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_40_DFFSR_129 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_9_DFFSR_27 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_7_AOI21X1_46 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_15_DFFSR_60 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_26_DFFSR_20 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_2_NAND3X1_175 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_3_DFFSR_205 INVX1_3/gnd DFFSR_79/S FILL
XFILL_2_BUFX2_95 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_30_DFFSR_132 INVX1_3/gnd DFFSR_79/S FILL
XFILL_24_5_1 AND2X2_38/B DFFSR_59/S FILL
XFILL_6_AOI21X1_49 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_44_DFFSR_236 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_7_DFFPOSX1_49 BUFX2_99/A DFFSR_92/S FILL
XFILL_20_DFFSR_135 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_6_4_0 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_5_AOI21X1_52 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_34_DFFSR_239 INVX1_39/gnd DFFSR_54/S FILL
XAOI21X1_49 AOI21X1_49/A AOI21X1_49/B BUFX2_36/Y BUFX2_7/gnd AOI21X1_49/Y DFFSR_216/S
+ AOI21X1
XFILL_10_DFFSR_138 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_4_AOI21X1_55 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_24_DFFSR_242 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_50_DFFSR_77 BUFX2_98/A DFFSR_32/S FILL
XFILL_3_NAND3X1_109 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_5_NOR2X1_14 INVX1_1/gnd DFFSR_97/S FILL
XFILL_4_6_1 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_3_AOI21X1_58 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_14_DFFSR_245 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_2_AOI21X1_61 AND2X2_38/B DFFSR_59/S FILL
XFILL_54_1 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_5_NAND2X1_145 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_34_DFFSR_27 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_6_DFFSR_74 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_6_DFFSR_132 INVX1_3/gnd DFFSR_79/S FILL
XFILL_1_AOI21X1_64 AND2X2_38/B DFFSR_59/S FILL
XFILL_23_DFFSR_67 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_47_DFFSR_163 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_0_AOI21X1_67 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_37_DFFSR_166 AND2X2_38/B DFFSR_59/S FILL
XBUFX2_52 BUFX2_53/A XOR2X1_1/gnd BUFX2_52/Y DFFSR_151/S BUFX2
XFILL_5_BUFX2_12 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_0_DFFSR_242 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_27_DFFSR_169 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_3_INVX1_216 INVX1_1/gnd DFFSR_97/S FILL
XFILL_41_DFFSR_273 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_17_DFFSR_172 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_31_DFFSR_276 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_9_AOI22X1_4 BUFX2_99/A DFFSR_92/S FILL
XFILL_1_NAND3X1_205 INVX1_1/gnd DFFSR_53/S FILL
XFILL_8_OAI21X1_91 BUFX2_8/gnd DFFSR_51/S FILL
XOAI21X1_2 INVX1_16/Y OAI21X1_4/B OAI21X1_2/C BUFX2_79/A OAI21X1_2/Y DFFSR_7/S OAI21X1
XFILL_7_OAI21X1_94 INVX1_67/gnd DFFSR_175/S FILL
XFILL_21_DFFSR_279 BUFX2_99/A DFFSR_7/S FILL
XFILL_3_INVX1_68 INVX1_67/gnd DFFSR_201/S FILL
XFILL_31_DFFSR_74 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_42_DFFSR_34 DFFSR_34/gnd DFFSR_34/S FILL
XNAND2X1_115 OAI22X1_52/Y NAND3X1_246/Y DFFSR_28/gnd NAND2X1_115/Y DFFSR_3/S NAND2X1
XFILL_3_XOR2X1_11 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_2_NOR2X1_51 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_6_OAI21X1_97 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_34_0_1 OR2X2_6/gnd DFFSR_53/S FILL
XOAI21X1_97 BUFX2_53/Y INVX1_194/Y OAI21X1_97/C BUFX2_72/gnd DFFSR_269/D DFFSR_276/S
+ OAI21X1
XFILL_15_DFFSR_24 BUFX2_98/A DFFSR_6/S FILL
XFILL_7_AOI21X1_10 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_2_NAND3X1_139 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_3_DFFSR_169 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_2_BUFX2_59 AND2X2_38/B DFFSR_23/S FILL
XFILL_6_AOI21X1_13 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_44_DFFSR_200 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_9_AND2X2_10 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_32_2_2 INVX1_1/gnd DFFSR_97/S FILL
XFILL_7_DFFSR_276 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_7_DFFPOSX1_13 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_5_AOI21X1_16 INVX1_67/gnd DFFSR_175/S FILL
XFILL_4_NAND2X1_175 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_6_NOR3X1_5 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_34_DFFSR_203 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_38_DFFSR_8 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_10_DFFSR_102 DFFSR_4/gnd DFFSR_98/S FILL
XAOI21X1_13 AOI21X1_13/A OAI21X1_41/Y AOI21X1_13/C DFFSR_34/gnd NOR3X1_5/C DFFSR_34/S
+ AOI21X1
XFILL_3_DFFPOSX1_2 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_4_AOI21X1_19 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_24_DFFSR_206 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_50_DFFSR_41 BUFX2_98/A DFFSR_6/S FILL
XFILL_39_DFFSR_81 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_2_DFFPOSX1_5 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_14_DFFSR_209 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_3_AOI21X1_22 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_16_DFFPOSX1_32 INVX1_67/gnd DFFSR_201/S FILL
XFILL_1_DFFPOSX1_8 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_2_AOI21X1_25 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_17_CLKBUF1_4 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_6_DFFSR_38 BUFX2_98/A DFFSR_6/S FILL
XFILL_23_DFFSR_31 BUFX2_79/A DFFSR_6/S FILL
XFILL_5_NAND2X1_109 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_12_DFFSR_71 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_1_AOI21X1_28 AND2X2_38/B DFFSR_23/S FILL
XFILL_0_NAND3X1_235 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_47_DFFSR_127 BUFX2_99/A DFFSR_92/S FILL
XFILL_0_AOI21X1_31 INVX1_39/gnd DFFSR_34/S FILL
XFILL_37_DFFSR_130 BUFX2_79/A DFFSR_6/S FILL
XFILL_0_DFFSR_206 OR2X2_2/gnd DFFSR_175/S FILL
XBUFX2_16 NOR2X1_7/Y BUFX2_98/A BUFX2_16/Y DFFSR_32/S BUFX2
XFILL_27_DFFSR_133 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_9_OAI21X1_52 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_16_XOR2X1_1 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_26_DFFPOSX1_21 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_3_INVX1_180 BUFX2_98/A DFFSR_6/S FILL
XFILL_41_DFFSR_237 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_47_DFFSR_88 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_3_CLKBUF1_1 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_17_DFFSR_136 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_8_OAI21X1_55 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_31_DFFSR_240 INVX1_39/gnd DFFSR_34/S FILL
XFILL_1_NAND3X1_169 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_21_DFFSR_243 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_6_NAND2X1_76 INVX1_3/gnd DFFSR_23/S FILL
XFILL_7_OAI21X1_58 INVX1_39/gnd DFFSR_54/S FILL
XFILL_3_INVX1_32 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_3_DFFSR_85 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_20_DFFSR_78 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_31_DFFSR_38 BUFX2_98/A DFFSR_6/S FILL
XFILL_6_DFFPOSX1_43 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_2_NOR2X1_15 BUFX2_99/A DFFSR_7/S FILL
XFILL_6_OAI21X1_61 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_5_NAND2X1_79 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_11_DFFSR_246 XOR2X1_1/gnd DFFSR_208/S FILL
XNAND2X1_76 BUFX2_57/Y AND2X2_33/B INVX1_3/gnd NAND2X1_77/B DFFSR_23/S NAND2X1
XFILL_5_OAI21X1_64 INVX1_1/gnd DFFSR_53/S FILL
XFILL_4_NAND2X1_82 DFFSR_1/gnd DFFSR_81/S FILL
XOAI21X1_61 OAI21X1_58/C OAI21X1_73/B AOI21X1_22/A DFFSR_1/gnd OAI21X1_61/Y DFFSR_1/S
+ OAI21X1
XFILL_3_DFFSR_133 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_3_NAND2X1_85 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_2_NAND3X1_103 AND2X2_38/B DFFSR_23/S FILL
XFILL_2_BUFX2_23 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_4_OAI21X1_67 INVX1_1/gnd DFFSR_97/S FILL
XFILL_44_DFFSR_164 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_3_OAI21X1_70 INVX1_3/gnd DFFSR_23/S FILL
XFILL_2_NAND2X1_88 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_7_DFFSR_240 INVX1_39/gnd DFFSR_34/S FILL
XFILL_14_XOR2X1_15 BUFX2_99/A DFFSR_7/S FILL
XFILL_4_NAND2X1_139 INVX1_1/gnd DFFSR_97/S FILL
XFILL_34_DFFSR_167 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_12_NOR3X1_2 INVX1_1/gnd DFFSR_53/S FILL
XFILL_1_NAND2X1_91 INVX1_39/gnd DFFSR_54/S FILL
XFILL_2_OAI21X1_73 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_48_DFFSR_271 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_24_DFFSR_170 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_0_NAND2X1_94 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_1_OAI21X1_76 INVX1_1/gnd DFFSR_53/S FILL
XFILL_38_DFFSR_274 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_39_DFFSR_45 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_0_INVX1_217 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_0_INVX1_79 INVX1_39/gnd DFFSR_54/S FILL
XFILL_28_DFFSR_85 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_14_DFFSR_173 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_28_DFFSR_277 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_0_OAI21X1_79 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_6_AOI22X1_5 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_18_DFFSR_280 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_12_DFFSR_35 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_0_XOR2X1_12 INVX1_3/gnd DFFSR_23/S FILL
XFILL_0_NAND3X1_199 INVX1_1/gnd DFFSR_97/S FILL
XFILL_0_DFFSR_170 OR2X2_6/gnd DFFSR_92/S FILL
XDFFSR_280 BUFX2_78/A DFFSR_79/CLK DFFSR_274/R DFFSR_53/S DFFSR_280/D OR2X2_6/gnd
+ DFFSR_53/S DFFSR
XFILL_25_DFFSR_2 BUFX2_79/A DFFSR_7/S FILL
XFILL_41_DFFSR_201 INVX1_67/gnd DFFSR_201/S FILL
XFILL_3_INVX1_144 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_47_DFFSR_52 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_6_AND2X2_11 BUFX2_99/A DFFSR_7/S FILL
XFILL_36_DFFSR_92 BUFX2_99/A DFFSR_92/S FILL
XFILL_17_DFFSR_100 INVX1_1/gnd DFFSR_97/S FILL
XFILL_4_DFFSR_277 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_8_OAI21X1_19 BUFX2_98/A DFFSR_32/S FILL
XFILL_31_DFFSR_204 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_1_NAND3X1_133 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_6_NAND2X1_40 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_7_OAI21X1_22 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_21_DFFSR_207 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_20_DFFSR_42 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_3_DFFSR_49 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_11_DFFSR_210 BUFX2_98/A DFFSR_6/S FILL
XFILL_3_NAND2X1_169 INVX1_1/gnd DFFSR_53/S FILL
XFILL_5_NAND2X1_43 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_6_OAI21X1_25 DFFSR_62/gnd DFFSR_62/S FILL
XNAND2X1_40 DFFSR_170/D AND2X2_18/Y OR2X2_6/gnd NAND3X1_76/A DFFSR_53/S NAND2X1
XFILL_5_OAI21X1_28 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_4_NAND2X1_46 INVX1_39/gnd DFFSR_34/S FILL
XFILL_14_CLKBUF1_5 BUFX2_99/A DFFSR_92/S FILL
XOAI21X1_25 XOR2X1_1/B NOR2X1_66/B OAI21X1_25/C DFFSR_62/gnd AOI21X1_7/A DFFSR_62/S
+ OAI21X1
XFILL_3_NAND2X1_49 INVX1_3/gnd DFFSR_79/S FILL
XFILL_4_OAI21X1_31 AND2X2_38/B DFFSR_23/S FILL
XDFFPOSX1_43 INVX1_133/A CLKBUF1_43/Y NOR2X1_77/Y OR2X2_2/gnd DFFSR_216/S DFFPOSX1
XFILL_44_DFFSR_128 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_3_OAI21X1_34 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_2_NAND2X1_52 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_44_DFFSR_99 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_15_DFFPOSX1_26 AND2X2_38/B DFFSR_23/S FILL
XFILL_7_DFFSR_204 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_4_NAND2X1_103 AND2X2_38/B DFFSR_23/S FILL
XFILL_34_DFFSR_131 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_2_OAI21X1_37 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_1_NAND2X1_55 INVX1_39/gnd DFFSR_34/S FILL
XFILL_48_DFFSR_235 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_24_DFFSR_134 INVX1_1/gnd DFFSR_53/S FILL
XFILL_5_AND2X2_8 BUFX2_99/A DFFSR_7/S FILL
XFILL_0_NAND2X1_58 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_1_OAI21X1_40 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_38_DFFSR_238 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_0_INVX1_43 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_0_DFFSR_96 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_0_INVX1_181 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_28_DFFSR_49 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_17_DFFSR_89 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_0_CLKBUF1_2 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_14_DFFSR_137 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_19_3 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_28_DFFSR_241 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_0_OAI21X1_43 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_9_XNOR2X1_4 BUFX2_98/A DFFSR_6/S FILL
XFILL_33_3_0 INVX1_1/gnd DFFSR_53/S FILL
XFILL_25_DFFPOSX1_15 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_18_DFFSR_244 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_0_NAND3X1_163 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_8_AOI22X1_12 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_31_5_1 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_7_AOI22X1_15 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_5_DFFPOSX1_37 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_0_DFFSR_134 INVX1_1/gnd DFFSR_53/S FILL
XDFFSR_244 INVX1_89/A CLKBUF1_17/Y BUFX2_69/Y DFFSR_81/S DFFSR_236/Q DFFSR_1/gnd DFFSR_81/S
+ DFFSR
XFILL_6_AOI22X1_18 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_41_DFFSR_165 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_3_INVX1_108 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_47_DFFSR_16 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_36_DFFSR_56 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_25_DFFSR_96 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_4_DFFSR_241 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_5_AOI22X1_21 AND2X2_38/B DFFSR_59/S FILL
XFILL_31_DFFSR_168 OR2X2_6/gnd DFFSR_92/S FILL
XAOI22X1_18 BUFX2_56/Y AND2X2_34/B INVX1_135/A INVX1_145/A OR2X2_1/gnd AOI22X1_18/Y
+ DFFSR_59/S AOI22X1
XFILL_45_DFFSR_272 INVX1_3/gnd DFFSR_23/S FILL
XFILL_4_AOI22X1_24 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_21_DFFSR_171 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_35_DFFSR_275 BUFX2_99/A DFFSR_92/S FILL
XFILL_3_DFFSR_13 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_3_AOI22X1_27 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_3_NAND2X1_133 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_11_DFFSR_174 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_3_AOI22X1_6 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_25_DFFSR_278 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_4_NAND2X1_10 BUFX2_79/A DFFSR_7/S FILL
XFILL_7_XOR2X1_10 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_6_NOR2X1_50 INVX1_39/gnd DFFSR_34/S FILL
XFILL_11_OAI22X1_51 INVX1_39/gnd DFFSR_54/S FILL
XFILL_3_NAND2X1_13 BUFX2_99/A DFFSR_92/S FILL
XFILL_44_DFFSR_63 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_2_NAND2X1_16 BUFX2_79/A DFFSR_7/S FILL
XFILL_7_DFFSR_168 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_1_OAI21X1_115 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_24_DFFPOSX1_45 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_1_NAND2X1_19 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_48_DFFSR_199 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_8_NAND3X1_75 BUFX2_79/A DFFSR_7/S FILL
XFILL_0_NAND2X1_22 BUFX2_99/A DFFSR_7/S FILL
XFILL_0_DFFSR_60 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_38_DFFSR_202 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_8_NAND3X1_248 INVX1_3/gnd DFFSR_79/S FILL
XFILL_0_INVX1_145 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_3_AND2X2_12 BUFX2_98/A DFFSR_32/S FILL
XFILL_28_DFFSR_13 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_17_DFFSR_53 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_14_DFFSR_101 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_7_NAND3X1_78 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_4_BUFX2_88 INVX1_3/gnd DFFSR_23/S FILL
XFILL_1_DFFSR_278 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_28_DFFSR_205 INVX1_3/gnd DFFSR_79/S FILL
XFILL_6_NAND3X1_81 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_18_DFFSR_208 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_41_0_1 BUFX2_98/A DFFSR_32/S FILL
XFILL_5_NAND3X1_84 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_0_NAND3X1_127 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_21_CLKBUF1_3 BUFX2_98/A DFFSR_6/S FILL
XNAND3X1_81 DFFSR_187/D BUFX2_29/Y BUFX2_25/Y DFFSR_1/gnd NAND3X1_84/B DFFSR_1/S NAND3X1
XFILL_9_NAND3X1_182 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_4_NAND3X1_87 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_16_DFFSR_9 BUFX2_79/A DFFSR_6/S FILL
XFILL_39_2_2 BUFX2_79/A DFFSR_6/S FILL
XFILL_11_CLKBUF1_6 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_51_DFFSR_126 BUFX2_99/A DFFSR_7/S FILL
XFILL_3_NAND3X1_90 OR2X2_1/gnd DFFSR_59/S FILL
XDFFSR_208 DFFSR_216/D CLKBUF1_14/Y BUFX2_64/Y DFFSR_208/S DFFSR_208/D DFFSR_62/gnd
+ DFFSR_208/S DFFSR
XFILL_2_NAND2X1_163 INVX1_67/gnd DFFSR_201/S FILL
XFILL_41_DFFSR_129 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_2_NAND3X1_93 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_25_DFFSR_60 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_36_DFFSR_20 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_8_DFFSR_67 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_4_DFFSR_205 INVX1_3/gnd DFFSR_79/S FILL
XFILL_31_DFFSR_132 INVX1_3/gnd DFFSR_79/S FILL
XFILL_1_NAND3X1_96 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_45_DFFSR_236 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_0_NAND3X1_99 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_21_DFFSR_135 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_14_DFFPOSX1_20 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_35_DFFSR_239 INVX1_39/gnd DFFSR_54/S FILL
XFILL_11_DFFSR_138 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_25_DFFSR_242 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_6_NOR2X1_14 INVX1_1/gnd DFFSR_97/S FILL
XFILL_24_8 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_37_DFFSR_5 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_15_DFFSR_245 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_10_OAI22X1_18 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_44_DFFSR_27 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_7_DFFSR_132 INVX1_3/gnd DFFSR_79/S FILL
XFILL_33_DFFSR_67 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_48_DFFSR_163 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_8_NAND3X1_39 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_9_OAI22X1_21 BUFX2_98/A DFFSR_32/S FILL
XFILL_0_INVX1_109 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_0_DFFSR_24 BUFX2_98/A DFFSR_6/S FILL
XFILL_38_DFFSR_166 AND2X2_38/B DFFSR_59/S FILL
XFILL_8_NAND3X1_212 INVX1_39/gnd DFFSR_54/S FILL
XFILL_17_DFFSR_17 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_7_NAND3X1_42 BUFX2_79/A DFFSR_6/S FILL
XFILL_4_BUFX2_52 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_1_DFFSR_242 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_8_OAI22X1_24 BUFX2_98/A DFFSR_32/S FILL
XFILL_4_DFFPOSX1_31 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_28_DFFSR_169 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_4_INVX1_216 INVX1_1/gnd DFFSR_97/S FILL
XFILL_42_DFFSR_273 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_7_OAI22X1_27 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_6_NAND3X1_45 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_18_DFFSR_172 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_32_DFFSR_276 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_5_NAND3X1_48 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_6_OAI22X1_30 OR2X2_6/gnd DFFSR_53/S FILL
XXOR2X1_14 XOR2X1_14/A XOR2X1_14/B INVX1_1/gnd XOR2X1_14/Y DFFSR_53/S XOR2X1
XNAND3X1_45 DFFSR_14/Q BUFX2_19/Y BUFX2_13/Y OR2X2_3/gnd NAND3X1_45/Y DFFSR_60/S NAND3X1
XFILL_22_DFFSR_279 BUFX2_99/A DFFSR_7/S FILL
XFILL_0_AOI22X1_7 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_4_NAND3X1_51 BUFX2_99/A DFFSR_7/S FILL
XFILL_5_OAI22X1_33 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_41_DFFSR_74 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_4_XOR2X1_11 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_3_NOR2X1_51 DFFSR_34/gnd DFFSR_34/S FILL
XOAI22X1_30 INVX1_73/Y OAI22X1_45/B INVX1_74/Y OAI22X1_45/D OR2X2_6/gnd NOR2X1_39/A
+ DFFSR_53/S OAI22X1
XFILL_13_DFFPOSX1_50 INVX1_1/gnd DFFSR_53/S FILL
XFILL_4_OAI22X1_36 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_3_NAND3X1_54 OR2X2_3/gnd DFFSR_60/S FILL
XDFFSR_172 DFFSR_172/Q DFFSR_1/CLK BUFX2_68/Y DFFSR_62/S DFFSR_164/Q DFFSR_46/gnd
+ DFFSR_62/S DFFSR
XFILL_2_NAND2X1_127 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_2_NAND3X1_57 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_3_OAI22X1_39 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_25_DFFSR_24 BUFX2_98/A DFFSR_6/S FILL
XFILL_8_DFFSR_31 BUFX2_79/A DFFSR_6/S FILL
XFILL_14_DFFSR_64 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_4_DFFSR_169 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_1_NAND3X1_60 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_1_BUFX2_99 BUFX2_99/A DFFSR_7/S FILL
XFILL_2_OAI22X1_42 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_45_DFFSR_200 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_0_NAND3X1_63 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_1_OAI22X1_45 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_8_DFFSR_276 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_0_OAI21X1_109 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_35_DFFSR_203 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_0_AND2X2_13 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_23_DFFPOSX1_39 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_11_DFFSR_102 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_0_OAI22X1_48 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_25_DFFSR_206 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_1_XOR2X1_1 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_49_DFFSR_81 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_15_DFFSR_209 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_7_NAND3X1_242 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_18_CLKBUF1_4 OR2X2_3/gnd DFFSR_60/S FILL
XINVX1_65 INVX1_65/A BUFX2_7/gnd INVX1_65/Y DFFSR_151/S INVX1
XFILL_5_DFFSR_78 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_33_DFFSR_31 BUFX2_79/A DFFSR_6/S FILL
XFILL_22_DFFSR_71 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_48_DFFSR_127 BUFX2_99/A DFFSR_92/S FILL
XFILL_13_0_2 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_38_DFFSR_130 BUFX2_79/A DFFSR_6/S FILL
XINVX1_183 DFFSR_3/D BUFX2_79/A INVX1_183/Y DFFSR_6/S INVX1
XFILL_8_NAND3X1_176 NOR3X1_6/gnd DFFSR_79/S FILL
XCLKBUF1_4 BUFX2_1/Y OR2X2_3/gnd CLKBUF1_4/Y DFFSR_60/S CLKBUF1
XFILL_1_DFFSR_206 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_4_BUFX2_16 BUFX2_98/A DFFSR_32/S FILL
XFILL_9_XOR2X1_8 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_28_DFFSR_133 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_1_NAND2X1_157 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_42_DFFSR_237 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_4_DFFSR_8 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_4_CLKBUF1_1 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_18_DFFSR_136 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_32_DFFSR_240 INVX1_39/gnd DFFSR_34/S FILL
XFILL_5_NAND3X1_12 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_22_DFFSR_243 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_4_NAND3X1_15 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_30_DFFSR_78 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_41_DFFSR_38 BUFX2_98/A DFFSR_6/S FILL
XFILL_2_INVX1_72 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_3_NOR2X1_15 BUFX2_99/A DFFSR_7/S FILL
XFILL_13_DFFPOSX1_14 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_12_DFFSR_246 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_3_NAND3X1_18 BUFX2_79/A DFFSR_7/S FILL
XDFFSR_136 DFFSR_136/Q CLKBUF1_27/Y BUFX2_61/Y DFFSR_79/S BUFX2_89/A NOR3X1_6/gnd
+ DFFSR_79/S DFFSR
XFILL_2_NAND3X1_21 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_14_DFFSR_28 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_4_DFFSR_133 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_1_BUFX2_63 BUFX2_98/A DFFSR_32/S FILL
XFILL_1_NAND3X1_24 INVX1_1/gnd DFFSR_97/S FILL
XFILL_45_DFFSR_164 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_0_NAND3X1_27 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_8_DFFSR_240 INVX1_39/gnd DFFSR_34/S FILL
XFILL_40_3_0 BUFX2_98/A DFFSR_6/S FILL
XFILL_15_XOR2X1_15 BUFX2_99/A DFFSR_7/S FILL
XFILL_35_DFFSR_167 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_49_DFFSR_271 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_0_OAI22X1_12 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_25_DFFSR_170 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_39_DFFSR_274 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_49_DFFSR_45 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_1_INVX1_217 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_38_DFFSR_85 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_38_5_1 BUFX2_79/A DFFSR_7/S FILL
XFILL_15_DFFSR_173 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_7_NAND3X1_206 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_29_DFFSR_277 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_7_AOI22X1_5 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_3_DFFPOSX1_25 BUFX2_79/A DFFSR_6/S FILL
XINVX1_29 DFFSR_28/Q DFFSR_28/gnd INVX1_29/Y DFFSR_8/S INVX1
XDFFSR_82 DFFSR_82/Q DFFSR_82/CLK DFFSR_35/R DFFSR_98/S INVX1_13/A BUFX2_77/gnd DFFSR_98/S
+ DFFSR
XFILL_5_DFFSR_42 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_19_DFFSR_280 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_22_DFFSR_35 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_11_DFFSR_75 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_1_XOR2X1_12 INVX1_3/gnd DFFSR_23/S FILL
XFILL_0_NOR2X1_52 DFFSR_1/gnd DFFSR_1/S FILL
XINVX1_147 INVX1_147/A BUFX2_7/gnd INVX1_147/Y DFFSR_216/S INVX1
XFILL_8_NAND3X1_140 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_1_DFFSR_170 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_12_DFFPOSX1_44 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_15_XOR2X1_5 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_42_DFFSR_201 INVX1_67/gnd DFFSR_201/S FILL
XFILL_49_DFFSR_8 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_1_NAND2X1_121 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_7_AND2X2_11 BUFX2_99/A DFFSR_7/S FILL
XFILL_46_DFFSR_92 BUFX2_99/A DFFSR_92/S FILL
XFILL_18_DFFSR_100 INVX1_1/gnd DFFSR_97/S FILL
XFILL_5_DFFSR_277 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_32_DFFSR_204 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_7_AND2X2_1 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_22_DFFSR_207 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_2_INVX1_36 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_30_DFFSR_42 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_2_DFFSR_89 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_19_DFFSR_82 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_12_DFFSR_210 BUFX2_98/A DFFSR_6/S FILL
XDFFSR_100 DFFSR_100/Q DFFSR_79/CLK DFFSR_7/R DFFSR_97/S DFFSR_92/Q INVX1_1/gnd DFFSR_97/S
+ DFFSR
XFILL_22_DFFPOSX1_33 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_15_CLKBUF1_5 BUFX2_99/A DFFSR_92/S FILL
XFILL_6_NAND3X1_236 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_1_BUFX2_27 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_45_DFFSR_128 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_8_DFFSR_204 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_35_DFFSR_131 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_11_NOR3X1_6 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_49_DFFSR_235 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_48_0_1 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_25_DFFSR_134 INVX1_1/gnd DFFSR_53/S FILL
XFILL_39_DFFSR_238 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_1_INVX1_181 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_38_DFFSR_49 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_27_DFFSR_89 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_1_CLKBUF1_2 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_15_DFFSR_137 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_7_NAND3X1_170 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_29_DFFSR_241 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_46_2_2 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_0_NAND2X1_151 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_19_DFFSR_244 DFFSR_1/gnd DFFSR_81/S FILL
XDFFSR_46 DFFSR_62/D AOI21X1_3/B DFFSR_1/R DFFSR_54/S DFFSR_46/D DFFSR_46/gnd DFFSR_54/S
+ DFFSR
XFILL_11_DFFSR_39 INVX1_3/gnd DFFSR_79/S FILL
XFILL_0_NOR2X1_16 BUFX2_79/A DFFSR_7/S FILL
XFILL_8_NAND3X1_104 AND2X2_38/B DFFSR_23/S FILL
XINVX1_111 DFFSR_144/D OR2X2_1/gnd INVX1_111/Y DFFSR_59/S INVX1
XFILL_1_DFFSR_134 INVX1_1/gnd DFFSR_53/S FILL
XFILL_15_DFFSR_6 BUFX2_79/A DFFSR_6/S FILL
XFILL_42_DFFSR_165 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_46_DFFSR_56 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_35_DFFSR_96 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_5_DFFSR_241 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_32_DFFSR_168 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_46_DFFSR_272 INVX1_3/gnd DFFSR_23/S FILL
XFILL_14_1_0 INVX1_39/gnd DFFSR_54/S FILL
XFILL_22_DFFSR_171 BUFX2_8/gnd DFFSR_81/S FILL
XAOI22X1_9 NOR3X1_4/Y DFFSR_225/Q DFFSR_217/Q NOR3X1_3/Y OR2X2_2/gnd AOI22X1_9/Y DFFSR_216/S
+ AOI22X1
XFILL_36_DFFSR_275 BUFX2_99/A DFFSR_92/S FILL
XFILL_2_DFFSR_53 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_19_DFFSR_46 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_6_BUFX2_81 BUFX2_79/A DFFSR_7/S FILL
XFILL_12_DFFSR_174 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_26_DFFSR_278 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_4_AOI22X1_6 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_12_3_1 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_8_XOR2X1_10 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_6_NAND3X1_200 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_20_CLKBUF1_36 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_10_5_2 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_19_CLKBUF1_39 INVX1_1/gnd DFFSR_53/S FILL
XFILL_36_DFFSR_2 BUFX2_79/A DFFSR_7/S FILL
XFILL_8_DFFSR_168 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_2_DFFPOSX1_19 DFFSR_34/gnd DFFSR_1/S FILL
XAND2X2_15 INVX1_63/Y NOR3X1_4/B INVX1_3/gnd AND2X2_15/Y DFFSR_23/S AND2X2
XFILL_18_CLKBUF1_42 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_49_DFFSR_199 XOR2X1_1/gnd DFFSR_208/S FILL
XNAND3X1_236 NAND3X1_233/Y NAND3X1_236/B OR2X2_3/Y DFFSR_4/gnd AOI21X1_37/A DFFSR_98/S
+ NAND3X1
XFILL_17_CLKBUF1_45 BUFX2_79/A DFFSR_7/S FILL
XFILL_39_DFFSR_202 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_1_INVX1_145 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_16_DFFSR_93 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_4_AND2X2_12 BUFX2_98/A DFFSR_32/S FILL
XFILL_38_DFFSR_13 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_27_DFFSR_53 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_15_DFFSR_101 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_7_NAND3X1_134 INVX1_39/gnd DFFSR_54/S FILL
XFILL_2_DFFSR_278 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_16_CLKBUF1_48 INVX1_3/gnd DFFSR_79/S FILL
XFILL_29_DFFSR_205 INVX1_3/gnd DFFSR_79/S FILL
XFILL_11_DFFPOSX1_38 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_0_NAND2X1_115 DFFSR_28/gnd DFFSR_3/S FILL
XDFFSR_10 DFFSR_66/D CLKBUF1_38/Y DFFSR_15/R DFFSR_5/S DFFSR_50/Q DFFSR_5/gnd DFFSR_5/S
+ DFFSR
XFILL_19_DFFSR_208 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_12_CLKBUF1_6 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_21_DFFPOSX1_27 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_42_DFFSR_129 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_35_DFFSR_60 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_46_DFFSR_20 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_5_DFFSR_205 INVX1_3/gnd DFFSR_79/S FILL
XFILL_32_DFFSR_132 INVX1_3/gnd DFFSR_79/S FILL
XFILL_5_NAND3X1_230 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_46_DFFSR_236 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_22_DFFSR_135 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_2_DFFSR_17 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_1_DFFPOSX1_49 BUFX2_99/A DFFSR_92/S FILL
XFILL_36_DFFSR_239 INVX1_39/gnd DFFSR_54/S FILL
XFILL_19_DFFSR_10 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_6_BUFX2_45 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_12_DFFSR_138 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_26_DFFSR_242 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_20_0_2 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_16_DFFSR_245 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_6_NAND3X1_164 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_8_DFFSR_132 INVX1_3/gnd DFFSR_79/S FILL
XFILL_43_DFFSR_67 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_49_DFFSR_163 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_0_1_2 BUFX2_72/gnd DFFSR_276/S FILL
XNAND3X1_200 INVX1_168/Y INVX1_167/Y OAI21X1_78/C OR2X2_6/gnd NAND3X1_201/A DFFSR_53/S
+ NAND3X1
XFILL_1_INVX1_109 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_39_DFFSR_166 AND2X2_38/B DFFSR_59/S FILL
XFILL_27_DFFSR_17 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_16_DFFSR_57 BUFX2_79/A DFFSR_6/S FILL
XFILL_3_BUFX2_92 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_2_DFFSR_242 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_16_CLKBUF1_12 AND2X2_38/B DFFSR_23/S FILL
XFILL_29_DFFSR_169 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_43_DFFSR_273 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_19_DFFSR_172 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_15_CLKBUF1_15 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_33_DFFSR_276 BUFX2_72/gnd DFFSR_276/S FILL
XNOR2X1_54 NOR2X1_54/A NOR2X1_54/B BUFX2_8/gnd NOR2X1_54/Y DFFSR_51/S NOR2X1
XFILL_14_CLKBUF1_18 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_3_DFFSR_5 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_1_AOI22X1_7 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_23_DFFSR_279 BUFX2_99/A DFFSR_7/S FILL
XFILL_13_CLKBUF1_21 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_5_XOR2X1_11 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_4_NOR2X1_51 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_47_3_0 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_12_CLKBUF1_24 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_7_OAI21X1_116 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_35_DFFSR_24 BUFX2_98/A DFFSR_6/S FILL
XFILL_7_DFFSR_71 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_24_DFFSR_64 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_11_CLKBUF1_27 INVX1_1/gnd DFFSR_97/S FILL
XFILL_5_DFFSR_169 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_45_5_1 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_10_CLKBUF1_30 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_46_DFFSR_200 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_5_NAND3X1_194 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_9_DFFSR_276 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_1_DFFPOSX1_13 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_1_OR2X2_5 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_36_DFFSR_203 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_1_AND2X2_13 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_12_DFFSR_102 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_26_DFFSR_206 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_9_CLKBUF1_33 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_16_DFFSR_209 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_27_DFFSR_9 BUFX2_79/A DFFSR_6/S FILL
XFILL_8_CLKBUF1_36 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_6_NAND3X1_128 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_7_CLKBUF1_39 INVX1_1/gnd DFFSR_53/S FILL
XFILL_10_DFFPOSX1_32 INVX1_67/gnd DFFSR_201/S FILL
XFILL_19_CLKBUF1_4 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_4_INVX1_65 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_43_DFFSR_31 BUFX2_79/A DFFSR_6/S FILL
XFILL_32_DFFSR_71 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_6_CLKBUF1_42 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_49_DFFSR_127 BUFX2_99/A DFFSR_92/S FILL
XFILL_5_CLKBUF1_45 BUFX2_79/A DFFSR_7/S FILL
XNAND3X1_164 INVX1_152/Y OAI21X1_46/C AOI21X1_20/B DFFSR_34/gnd AOI21X1_13/A DFFSR_1/S
+ NAND3X1
XFILL_39_DFFSR_130 BUFX2_79/A DFFSR_6/S FILL
XCLKBUF1_42 BUFX2_2/Y DFFSR_4/gnd DFFSR_45/CLK DFFSR_98/S CLKBUF1
XFILL_16_DFFSR_21 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_4_CLKBUF1_48 INVX1_3/gnd DFFSR_79/S FILL
XFILL_2_DFFSR_206 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_3_BUFX2_56 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_29_DFFSR_133 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_11_6_0 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_43_DFFSR_237 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_20_DFFPOSX1_21 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_5_CLKBUF1_1 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_19_DFFSR_136 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_7_NOR3X1_2 INVX1_1/gnd DFFSR_53/S FILL
XFILL_33_DFFSR_240 INVX1_39/gnd DFFSR_34/S FILL
XNOR2X1_18 NOR2X1_18/A NOR2X1_18/B OR2X2_4/gnd NOR2X1_18/Y DFFSR_3/S NOR2X1
XFILL_48_DFFSR_5 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_23_DFFSR_243 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_4_NAND3X1_224 INVX1_39/gnd DFFSR_54/S FILL
XFILL_40_DFFSR_78 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_4_NOR2X1_15 BUFX2_99/A DFFSR_7/S FILL
XFILL_0_DFFPOSX1_43 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_13_DFFSR_246 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_7_DFFSR_35 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_50_5 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_24_DFFSR_28 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_5_DFFSR_133 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_13_DFFSR_68 BUFX2_98/A DFFSR_6/S FILL
XFILL_46_DFFSR_164 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_5_NAND3X1_158 AND2X2_38/B DFFSR_59/S FILL
XFILL_53_2_2 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_9_DFFSR_240 INVX1_39/gnd DFFSR_34/S FILL
XFILL_36_DFFSR_167 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_3_INVX1_7 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_50_DFFSR_271 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_0_XOR2X1_5 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_26_DFFSR_170 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_40_DFFSR_274 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_48_DFFSR_85 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_2_INVX1_217 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_16_DFFSR_173 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_30_DFFSR_277 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_8_AOI22X1_5 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_20_DFFSR_280 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_32_DFFSR_35 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_4_INVX1_29 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_4_DFFSR_82 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_21_DFFSR_75 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_2_XOR2X1_12 INVX1_3/gnd DFFSR_23/S FILL
XFILL_1_NOR2X1_52 DFFSR_1/gnd DFFSR_1/S FILL
XNAND3X1_128 NOR2X1_56/Y NOR2X1_57/Y NOR2X1_58/Y NOR3X1_6/gnd XNOR2X1_4/B DFFSR_79/S
+ NAND3X1
XFILL_21_1_0 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_4_CLKBUF1_12 AND2X2_38/B DFFSR_23/S FILL
XFILL_3_BUFX2_20 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_2_DFFSR_170 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_43_DFFSR_201 INVX1_67/gnd DFFSR_201/S FILL
XFILL_3_CLKBUF1_15 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_8_AND2X2_11 BUFX2_99/A DFFSR_7/S FILL
XFILL_19_DFFSR_100 INVX1_1/gnd DFFSR_97/S FILL
XFILL_19_3_1 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_6_DFFSR_277 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_6_OAI21X1_110 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_33_DFFSR_204 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_14_DFFSR_3 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_2_CLKBUF1_18 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_1_2_0 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_4_NAND3X1_188 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_1_CLKBUF1_21 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_23_DFFSR_207 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_40_DFFSR_42 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_1_INVX1_76 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_29_DFFSR_82 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_17_5_2 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_0_CLKBUF1_24 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_13_DFFSR_210 BUFX2_98/A DFFSR_6/S FILL
XFILL_16_CLKBUF1_5 BUFX2_99/A DFFSR_92/S FILL
XFILL_13_DFFSR_32 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_0_BUFX2_67 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_5_NAND3X1_122 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_46_DFFSR_128 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_9_DFFSR_204 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_36_DFFSR_131 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_50_DFFSR_235 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_26_DFFSR_134 INVX1_1/gnd DFFSR_53/S FILL
XFILL_10_2 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_40_DFFSR_238 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_48_DFFSR_49 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_37_DFFSR_89 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_2_INVX1_181 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_2_CLKBUF1_2 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_16_DFFSR_137 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_30_DFFSR_241 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_20_DFFSR_244 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_21_DFFSR_39 INVX1_3/gnd DFFSR_79/S FILL
XFILL_4_DFFSR_46 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_19_DFFPOSX1_15 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_1_NOR2X1_16 BUFX2_79/A DFFSR_7/S FILL
XFILL_10_DFFSR_79 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_10_DFFSR_247 BUFX2_99/A DFFSR_7/S FILL
XFILL_3_NAND3X1_218 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_2_DFFSR_134 INVX1_1/gnd DFFSR_53/S FILL
XFILL_27_DFFPOSX1_3 INVX1_39/gnd DFFSR_34/S FILL
XFILL_43_DFFSR_165 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_14_XOR2X1_9 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_45_DFFSR_96 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_6_DFFSR_241 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_26_DFFPOSX1_6 AND2X2_38/B DFFSR_23/S FILL
XFILL_33_DFFSR_168 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_27_0_2 INVX1_3/gnd DFFSR_79/S FILL
XFILL_47_DFFSR_272 INVX1_3/gnd DFFSR_23/S FILL
XFILL_25_DFFPOSX1_9 INVX1_67/gnd DFFSR_201/S FILL
XFILL_23_DFFSR_171 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_6_AND2X2_5 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_4_NAND3X1_152 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_1_INVX1_40 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_37_DFFSR_275 BUFX2_99/A DFFSR_92/S FILL
XFILL_1_DFFSR_93 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_18_DFFSR_86 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_29_DFFSR_46 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_13_DFFSR_174 BUFX2_8/gnd DFFSR_51/S FILL
XOAI21X1_110 NOR3X1_6/B NOR3X1_6/C INVX1_209/Y NOR3X1_6/gnd AOI21X1_63/C DFFSR_91/S
+ OAI21X1
XFILL_5_AOI22X1_6 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_9_DFFPOSX1_26 AND2X2_38/B DFFSR_23/S FILL
XFILL_27_DFFSR_278 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_9_XOR2X1_10 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_7_1_2 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_0_BUFX2_31 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_0_OAI21X1_1 BUFX2_79/A DFFSR_7/S FILL
XFILL_9_DFFSR_168 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_18_DFFPOSX1_45 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_50_DFFSR_199 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_40_DFFSR_202 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_2_INVX1_145 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_26_DFFSR_93 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_5_AND2X2_12 BUFX2_98/A DFFSR_32/S FILL
XFILL_48_DFFSR_13 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_37_DFFSR_53 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_16_DFFSR_101 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_2_NAND3X1_248 INVX1_3/gnd DFFSR_79/S FILL
XFILL_3_DFFSR_278 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_30_DFFSR_205 INVX1_3/gnd DFFSR_79/S FILL
XFILL_54_3_0 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_20_DFFSR_208 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_4_DFFSR_10 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_5_OAI21X1_104 INVX1_67/gnd DFFSR_201/S FILL
XFILL_10_DFFSR_43 BUFX2_98/A DFFSR_6/S FILL
XFILL_10_DFFSR_211 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_52_5_1 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_3_NAND3X1_182 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_13_CLKBUF1_6 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_2_DFFSR_2 BUFX2_79/A DFFSR_7/S FILL
XFILL_43_DFFSR_129 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_45_DFFSR_60 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_6_DFFSR_205 INVX1_3/gnd DFFSR_79/S FILL
XFILL_33_DFFSR_132 INVX1_3/gnd DFFSR_79/S FILL
XFILL_47_DFFSR_236 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_23_DFFSR_135 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_4_NAND3X1_116 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_1_DFFSR_57 BUFX2_79/A DFFSR_6/S FILL
XFILL_37_DFFSR_239 INVX1_39/gnd DFFSR_54/S FILL
XFILL_29_DFFSR_10 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_18_DFFSR_50 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_5_BUFX2_85 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_13_DFFSR_138 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_27_DFFSR_242 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_32_2 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_0_OR2X2_2 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_6_NAND2X1_152 INVX1_1/gnd DFFSR_97/S FILL
XFILL_17_DFFSR_245 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_26_DFFSR_6 BUFX2_79/A DFFSR_6/S FILL
XFILL_9_DFFSR_132 INVX1_3/gnd DFFSR_79/S FILL
XFILL_18_6_0 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_50_DFFSR_163 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_2_INVX1_109 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_40_DFFSR_166 AND2X2_38/B DFFSR_59/S FILL
XFILL_37_DFFSR_17 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_9_DFFSR_64 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_26_DFFSR_57 BUFX2_79/A DFFSR_6/S FILL
XFILL_15_DFFSR_97 INVX1_1/gnd DFFSR_97/S FILL
XFILL_2_NAND3X1_212 INVX1_39/gnd DFFSR_54/S FILL
XFILL_3_DFFSR_242 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_30_DFFSR_169 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_44_DFFSR_273 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_20_DFFSR_172 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_34_DFFSR_276 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_10_DFFSR_175 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_2_AOI22X1_7 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_24_DFFSR_279 BUFX2_99/A DFFSR_7/S FILL
XFILL_15_DFFPOSX1_3 INVX1_39/gnd DFFSR_34/S FILL
XFILL_6_XOR2X1_11 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_3_NAND3X1_146 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_5_NOR2X1_51 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_47_DFFSR_2 BUFX2_79/A DFFSR_7/S FILL
XFILL_14_DFFPOSX1_6 AND2X2_38/B DFFSR_23/S FILL
XFILL_13_DFFPOSX1_9 INVX1_67/gnd DFFSR_201/S FILL
XFILL_8_DFFPOSX1_20 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_5_NAND2X1_182 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_34_DFFSR_64 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_45_DFFSR_24 BUFX2_98/A DFFSR_6/S FILL
XFILL_6_DFFSR_169 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_47_DFFSR_200 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_1_DFFSR_21 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_37_DFFSR_203 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_18_DFFSR_14 INVX1_1/gnd DFFSR_53/S FILL
XFILL_2_AND2X2_13 DFFSR_28/gnd DFFSR_3/S FILL
XBUFX2_89 BUFX2_89/A INVX1_1/gnd BUFX2_89/Y DFFSR_97/S BUFX2
XFILL_13_DFFSR_102 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_0_DFFSR_279 BUFX2_99/A DFFSR_7/S FILL
XFILL_5_BUFX2_49 INVX1_1/gnd DFFSR_97/S FILL
XFILL_17_DFFPOSX1_39 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_27_DFFSR_206 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_6_NAND2X1_116 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_2_INVX1_4 BUFX2_99/A DFFSR_7/S FILL
XFILL_17_DFFSR_209 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_28_1_0 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_1_NAND3X1_242 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_0_NOR2X1_2 INVX1_1/gnd DFFSR_97/S FILL
XFILL_42_DFFSR_71 XOR2X1_4/gnd DFFSR_91/S FILL
XNAND2X1_152 NAND2X1_151/B INVX1_208/Y INVX1_1/gnd AOI21X1_52/A DFFSR_97/S NAND2X1
XFILL_10_CLKBUF1_7 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_26_3_1 INVX1_3/gnd DFFSR_23/S FILL
XFILL_50_DFFSR_127 BUFX2_99/A DFFSR_92/S FILL
XFILL_27_DFFPOSX1_28 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_8_AOI21X1_44 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_40_DFFSR_130 BUFX2_79/A DFFSR_6/S FILL
XFILL_7_AOI21X1_47 INVX1_67/gnd DFFSR_175/S FILL
XFILL_8_2_0 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_9_DFFSR_28 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_26_DFFSR_21 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_15_DFFSR_61 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_2_NAND3X1_176 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_3_DFFSR_206 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_30_DFFSR_133 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_2_BUFX2_96 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_24_5_2 AND2X2_38/B DFFSR_59/S FILL
XFILL_6_AOI21X1_50 INVX1_67/gnd DFFSR_175/S FILL
XFILL_44_DFFSR_237 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_6_CLKBUF1_1 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_7_DFFPOSX1_50 INVX1_1/gnd DFFSR_53/S FILL
XFILL_20_DFFSR_136 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_6_4_1 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_5_AOI21X1_53 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_34_DFFSR_240 INVX1_39/gnd DFFSR_34/S FILL
XAOI21X1_50 AOI21X1_50/A AOI21X1_50/B BUFX2_36/Y INVX1_67/gnd AOI21X1_50/Y DFFSR_175/S
+ AOI21X1
XFILL_10_DFFSR_139 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_4_AOI21X1_56 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_24_DFFSR_243 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_3_NAND3X1_110 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_50_DFFSR_78 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_5_NOR2X1_15 BUFX2_99/A DFFSR_7/S FILL
XFILL_3_AOI21X1_59 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_4_6_2 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_14_DFFSR_246 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_2_AOI21X1_62 INVX1_3/gnd DFFSR_23/S FILL
XFILL_54_2 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_5_NAND2X1_146 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_34_DFFSR_28 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_23_DFFSR_68 BUFX2_98/A DFFSR_6/S FILL
XFILL_6_DFFSR_75 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_6_DFFSR_133 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_1_AOI21X1_65 INVX1_3/gnd DFFSR_23/S FILL
XFILL_47_DFFSR_164 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_0_AOI21X1_68 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_37_DFFSR_167 OR2X2_2/gnd DFFSR_216/S FILL
XBUFX2_53 BUFX2_53/A BUFX2_7/gnd BUFX2_53/Y DFFSR_216/S BUFX2
XFILL_51_DFFSR_271 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_0_DFFSR_243 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_5_BUFX2_13 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_27_DFFSR_170 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_41_DFFSR_274 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_3_INVX1_217 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_17_DFFSR_173 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_8_OAI21X1_92 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_31_DFFSR_277 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_9_AOI22X1_5 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_1_NAND3X1_206 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_7_OAI21X1_95 BUFX2_7/gnd DFFSR_216/S FILL
XOAI21X1_3 INVX1_23/Y OAI21X1_4/B OAI21X1_3/C BUFX2_99/A NOR2X1_13/B DFFSR_92/S OAI21X1
XFILL_21_DFFSR_280 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_42_DFFSR_35 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_3_INVX1_69 INVX1_3/gnd DFFSR_23/S FILL
XFILL_3_XOR2X1_12 INVX1_3/gnd DFFSR_23/S FILL
XFILL_31_DFFSR_75 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_2_NOR2X1_52 DFFSR_1/gnd DFFSR_1/S FILL
XNAND2X1_116 din[0] DFFSR_54/S DFFSR_46/gnd OAI21X1_85/C DFFSR_62/S NAND2X1
XFILL_6_OAI21X1_98 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_34_0_2 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_7_AOI21X1_11 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_15_DFFSR_25 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_2_NAND3X1_140 DFFSR_1/gnd DFFSR_1/S FILL
XOAI21X1_98 BUFX2_52/Y INVX1_195/Y OAI21X1_98/C DFFSR_46/gnd DFFSR_270/D DFFSR_54/S
+ OAI21X1
XFILL_3_DFFSR_170 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_2_BUFX2_60 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_6_AOI21X1_14 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_44_DFFSR_201 INVX1_67/gnd DFFSR_201/S FILL
XFILL_20_DFFSR_100 INVX1_1/gnd DFFSR_97/S FILL
XFILL_7_DFFSR_277 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_7_DFFPOSX1_14 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_34_DFFSR_204 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_5_AOI21X1_17 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_4_NAND2X1_176 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_6_NOR3X1_6 NOR3X1_6/gnd DFFSR_79/S FILL
XAOI21X1_14 AOI21X1_14/A AOI21X1_14/B AOI21X1_8/Y BUFX2_8/gnd AOI21X1_15/C DFFSR_81/S
+ AOI21X1
XFILL_10_DFFSR_103 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_38_DFFSR_9 BUFX2_79/A DFFSR_6/S FILL
XFILL_4_AOI21X1_20 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_3_DFFPOSX1_3 INVX1_39/gnd DFFSR_34/S FILL
XFILL_24_DFFSR_207 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_39_DFFSR_82 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_50_DFFSR_42 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_2_DFFPOSX1_6 AND2X2_38/B DFFSR_23/S FILL
XFILL_3_AOI21X1_23 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_14_DFFSR_210 BUFX2_98/A DFFSR_6/S FILL
XFILL_1_DFFPOSX1_9 INVX1_67/gnd DFFSR_201/S FILL
XFILL_16_DFFPOSX1_33 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_2_AOI21X1_26 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_17_CLKBUF1_5 BUFX2_99/A DFFSR_92/S FILL
XFILL_5_NAND2X1_110 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_6_DFFSR_39 INVX1_3/gnd DFFSR_79/S FILL
XFILL_12_DFFSR_72 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_23_DFFSR_32 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_1_AOI21X1_29 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_0_NAND3X1_236 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_47_DFFSR_128 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_0_AOI21X1_32 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_37_DFFSR_131 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_51_DFFSR_235 OR2X2_2/gnd DFFSR_216/S FILL
XBUFX2_17 NOR2X1_7/Y DFFSR_8/gnd BUFX2_17/Y DFFSR_8/S BUFX2
XFILL_0_DFFSR_207 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_27_DFFSR_134 INVX1_1/gnd DFFSR_53/S FILL
XFILL_41_DFFSR_238 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_26_DFFPOSX1_22 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_47_DFFSR_89 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_3_INVX1_181 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_3_CLKBUF1_2 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_17_DFFSR_137 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_8_OAI21X1_56 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_31_DFFSR_241 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_1_NAND3X1_170 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_6_NAND2X1_77 AND2X2_38/B DFFSR_23/S FILL
XFILL_7_OAI21X1_59 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_21_DFFSR_244 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_3_INVX1_33 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_3_DFFSR_86 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_31_DFFSR_39 INVX1_3/gnd DFFSR_79/S FILL
XFILL_6_DFFPOSX1_44 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_20_DFFSR_79 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_2_NOR2X1_16 BUFX2_79/A DFFSR_7/S FILL
XFILL_5_NAND2X1_80 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_11_DFFSR_247 BUFX2_99/A DFFSR_7/S FILL
XFILL_6_OAI21X1_62 INVX1_3/gnd DFFSR_79/S FILL
XNAND2X1_77 NAND2X1_77/A NAND2X1_77/B AND2X2_38/B AOI22X1_21/C DFFSR_23/S NAND2X1
XFILL_5_OAI21X1_65 INVX1_1/gnd DFFSR_53/S FILL
XFILL_4_NAND2X1_83 DFFSR_34/gnd DFFSR_34/S FILL
XOAI21X1_62 INVX1_146/Y INVX1_159/Y XOR2X1_4/A INVX1_3/gnd OAI21X1_62/Y DFFSR_79/S
+ OAI21X1
XFILL_2_NAND3X1_104 AND2X2_38/B DFFSR_23/S FILL
XFILL_4_OAI21X1_68 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_3_DFFSR_134 INVX1_1/gnd DFFSR_53/S FILL
XFILL_3_NAND2X1_86 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_2_BUFX2_24 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_44_DFFSR_165 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_3_OAI21X1_71 INVX1_3/gnd DFFSR_79/S FILL
XFILL_2_NAND2X1_89 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_7_DFFSR_241 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_4_NAND2X1_140 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_34_DFFSR_168 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_12_NOR3X1_3 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_1_NAND2X1_92 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_48_DFFSR_272 INVX1_3/gnd DFFSR_23/S FILL
XFILL_2_OAI21X1_74 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_24_DFFSR_171 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_1_OAI21X1_77 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_0_NAND2X1_95 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_28_DFFSR_86 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_38_DFFSR_275 BUFX2_99/A DFFSR_92/S FILL
XFILL_0_INVX1_80 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_39_DFFSR_46 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_25_6_0 AND2X2_38/B DFFSR_23/S FILL
XFILL_14_DFFSR_174 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_0_OAI21X1_80 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_6_AOI22X1_6 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_28_DFFSR_278 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_12_DFFSR_36 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_0_XOR2X1_13 INVX1_1/gnd DFFSR_97/S FILL
XFILL_1_OAI21X1_1 BUFX2_79/A DFFSR_7/S FILL
XFILL_0_NAND3X1_200 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_51_DFFSR_199 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_0_DFFSR_171 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_25_DFFSR_3 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_41_DFFSR_202 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_47_DFFSR_53 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_3_INVX1_145 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_36_DFFSR_93 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_6_AND2X2_12 BUFX2_98/A DFFSR_32/S FILL
XFILL_17_DFFSR_101 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_4_DFFSR_278 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_8_OAI21X1_20 AND2X2_38/B DFFSR_23/S FILL
XFILL_31_DFFSR_205 INVX1_3/gnd DFFSR_79/S FILL
XFILL_1_NAND3X1_134 INVX1_39/gnd DFFSR_54/S FILL
XFILL_7_OAI21X1_23 INVX1_67/gnd DFFSR_201/S FILL
XFILL_6_NAND2X1_41 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_21_DFFSR_208 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_3_DFFSR_50 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_20_DFFSR_43 BUFX2_98/A DFFSR_6/S FILL
XFILL_5_NAND2X1_44 INVX1_39/gnd DFFSR_34/S FILL
XFILL_6_OAI21X1_26 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_11_DFFSR_211 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_3_NAND2X1_170 BUFX2_7/gnd DFFSR_216/S FILL
XNAND2X1_41 DFFSR_235/Q NOR2X1_34/Y BUFX2_7/gnd NAND2X1_41/Y DFFSR_151/S NAND2X1
XFILL_5_OAI21X1_29 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_4_NAND2X1_47 DFFSR_62/gnd DFFSR_208/S FILL
XOAI21X1_26 XOR2X1_2/B XOR2X1_2/A OAI21X1_26/C OR2X2_2/gnd INVX1_140/A DFFSR_175/S
+ OAI21X1
XFILL_14_CLKBUF1_6 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_4_OAI21X1_32 AND2X2_38/B DFFSR_59/S FILL
XFILL_3_NAND2X1_50 DFFSR_62/gnd DFFSR_62/S FILL
XDFFPOSX1_44 AND2X2_35/A CLKBUF1_47/Y INVX1_213/Y OR2X2_2/gnd DFFSR_216/S DFFPOSX1
XFILL_44_DFFSR_129 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_3_OAI21X1_35 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_15_DFFPOSX1_27 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_2_NAND2X1_53 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_7_DFFSR_205 INVX1_3/gnd DFFSR_79/S FILL
XFILL_4_NAND2X1_104 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_34_DFFSR_132 INVX1_3/gnd DFFSR_79/S FILL
XFILL_1_NAND2X1_56 AND2X2_38/B DFFSR_59/S FILL
XFILL_2_OAI21X1_38 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_48_DFFSR_236 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_35_1_0 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_5_AND2X2_9 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_24_DFFSR_135 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_1_OAI21X1_41 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_38_DFFSR_239 INVX1_39/gnd DFFSR_54/S FILL
XFILL_0_NAND2X1_59 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_39_DFFSR_10 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_0_INVX1_182 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_28_DFFSR_50 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_0_INVX1_44 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_0_DFFSR_97 INVX1_1/gnd DFFSR_97/S FILL
XFILL_17_DFFSR_90 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_0_CLKBUF1_3 BUFX2_98/A DFFSR_6/S FILL
XFILL_14_DFFSR_138 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_19_4 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_0_OAI21X1_44 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_28_DFFSR_242 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_33_3_1 INVX1_1/gnd DFFSR_53/S FILL
XFILL_25_DFFPOSX1_16 INVX1_67/gnd DFFSR_175/S FILL
XFILL_18_DFFSR_245 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_9_AOI22X1_10 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_1_INVX1_1 INVX1_1/gnd DFFSR_53/S FILL
XFILL_8_AOI22X1_13 AND2X2_38/B DFFSR_23/S FILL
XFILL_0_NAND3X1_164 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_31_5_2 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_7_AOI22X1_16 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_5_DFFPOSX1_38 OR2X2_1/gnd DFFSR_51/S FILL
XDFFSR_245 INVX1_96/A CLKBUF1_6/Y BUFX2_66/Y DFFSR_34/S DFFSR_245/D DFFSR_34/gnd DFFSR_34/S
+ DFFSR
XFILL_0_DFFSR_135 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_6_AOI22X1_19 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_41_DFFSR_166 AND2X2_38/B DFFSR_59/S FILL
XFILL_47_DFFSR_17 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_3_INVX1_109 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_36_DFFSR_57 BUFX2_79/A DFFSR_6/S FILL
XFILL_25_DFFSR_97 INVX1_1/gnd DFFSR_97/S FILL
XFILL_4_DFFSR_242 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_5_AOI22X1_22 INVX1_3/gnd DFFSR_79/S FILL
XFILL_31_DFFSR_169 DFFSR_62/gnd DFFSR_62/S FILL
XAOI22X1_19 AND2X2_29/Y AND2X2_34/Y AOI22X1_19/C INVX1_144/Y OR2X2_1/gnd AOI21X1_10/C
+ DFFSR_51/S AOI22X1
XFILL_45_DFFSR_273 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_4_AOI22X1_25 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_21_DFFSR_172 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_3_DFFSR_14 INVX1_1/gnd DFFSR_53/S FILL
XFILL_35_DFFSR_276 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_3_AOI22X1_28 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_11_DFFSR_175 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_3_NAND2X1_134 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_3_AOI22X1_7 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_25_DFFSR_279 BUFX2_99/A DFFSR_7/S FILL
XFILL_4_NAND2X1_11 BUFX2_98/A DFFSR_6/S FILL
XFILL_7_XOR2X1_11 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_6_NOR2X1_51 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_3_NAND2X1_14 BUFX2_98/A DFFSR_32/S FILL
XFILL_2_NAND2X1_17 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_44_DFFSR_64 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_1_OAI21X1_116 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_7_DFFSR_169 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_24_DFFPOSX1_46 INVX1_39/gnd DFFSR_34/S FILL
XFILL_1_NAND2X1_20 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_9_NAND3X1_73 INVX1_1/gnd DFFSR_97/S FILL
XFILL_48_DFFSR_200 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_8_NAND3X1_76 INVX1_1/gnd DFFSR_53/S FILL
XFILL_0_NAND2X1_23 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_38_DFFSR_203 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_0_DFFSR_61 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_8_NAND3X1_249 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_28_DFFSR_14 INVX1_1/gnd DFFSR_53/S FILL
XFILL_0_INVX1_146 INVX1_3/gnd DFFSR_79/S FILL
XFILL_17_DFFSR_54 INVX1_39/gnd DFFSR_54/S FILL
XFILL_3_AND2X2_13 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_14_DFFSR_102 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_1_DFFSR_279 BUFX2_99/A DFFSR_7/S FILL
XFILL_7_NAND3X1_79 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_4_BUFX2_89 INVX1_1/gnd DFFSR_97/S FILL
XFILL_28_DFFSR_206 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_6_NAND3X1_82 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_18_DFFSR_209 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_41_0_2 BUFX2_98/A DFFSR_32/S FILL
XFILL_5_NAND3X1_85 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_0_NAND3X1_128 NOR3X1_6/gnd DFFSR_79/S FILL
XNAND3X1_82 DFFSR_155/D AND2X2_18/B BUFX2_28/Y DFFSR_1/gnd AND2X2_21/B DFFSR_1/S NAND3X1
XFILL_4_NAND3X1_88 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_11_CLKBUF1_7 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_3_NAND3X1_91 AND2X2_38/B DFFSR_59/S FILL
XDFFSR_209 INVX1_64/A CLKBUF1_34/Y BUFX2_62/Y DFFSR_276/S INVX1_65/A BUFX2_72/gnd
+ DFFSR_276/S DFFSR
XFILL_2_NAND2X1_164 INVX1_67/gnd DFFSR_175/S FILL
XFILL_41_DFFSR_130 BUFX2_79/A DFFSR_6/S FILL
XFILL_8_DFFSR_68 BUFX2_98/A DFFSR_6/S FILL
XFILL_2_NAND3X1_94 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_25_DFFSR_61 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_36_DFFSR_21 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_4_DFFSR_206 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_31_DFFSR_133 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_1_NAND3X1_97 AND2X2_38/B DFFSR_59/S FILL
XFILL_45_DFFSR_237 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_7_CLKBUF1_1 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_21_DFFSR_136 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_14_DFFPOSX1_21 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_35_DFFSR_240 INVX1_39/gnd DFFSR_34/S FILL
XFILL_11_DFFSR_139 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_25_DFFSR_243 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_6_NOR2X1_15 BUFX2_99/A DFFSR_7/S FILL
XFILL_24_9 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_15_DFFSR_246 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_37_DFFSR_6 BUFX2_79/A DFFSR_6/S FILL
XFILL_11_OAI22X1_16 AND2X2_38/B DFFSR_59/S FILL
XFILL_10_OAI22X1_19 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_44_DFFSR_28 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_33_DFFSR_68 BUFX2_98/A DFFSR_6/S FILL
XFILL_7_DFFSR_133 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_24_DFFPOSX1_10 INVX1_67/gnd DFFSR_201/S FILL
XFILL_48_DFFSR_164 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_9_OAI22X1_22 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_8_NAND3X1_40 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_38_DFFSR_167 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_0_DFFSR_25 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_0_INVX1_110 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_17_DFFSR_18 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_8_NAND3X1_213 INVX1_39/gnd DFFSR_54/S FILL
XFILL_1_DFFSR_243 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_7_NAND3X1_43 BUFX2_99/A DFFSR_7/S FILL
XFILL_8_OAI22X1_25 INVX1_39/gnd DFFSR_54/S FILL
XFILL_4_BUFX2_53 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_4_DFFPOSX1_32 INVX1_67/gnd DFFSR_201/S FILL
XFILL_28_DFFSR_170 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_42_DFFSR_274 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_6_NAND3X1_46 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_7_OAI22X1_28 INVX1_3/gnd DFFSR_23/S FILL
XFILL_18_DFFSR_173 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_32_DFFSR_277 BUFX2_72/gnd DFFSR_201/S FILL
XXOR2X1_15 XOR2X1_15/A XOR2X1_15/B BUFX2_99/A XOR2X1_15/Y DFFSR_7/S XOR2X1
XFILL_5_NAND3X1_49 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_6_OAI22X1_31 DFFSR_1/gnd DFFSR_81/S FILL
XNAND3X1_46 DFFSR_70/Q BUFX2_15/Y NOR2X1_2/Y DFFSR_4/gnd NAND3X1_47/B DFFSR_4/S NAND3X1
XFILL_0_AOI22X1_8 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_22_DFFSR_280 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_4_NAND3X1_52 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_5_OAI22X1_34 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_4_XOR2X1_12 INVX1_3/gnd DFFSR_23/S FILL
XFILL_41_DFFSR_75 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_3_NOR2X1_52 DFFSR_1/gnd DFFSR_1/S FILL
XOAI22X1_31 INVX1_76/Y OAI22X1_43/B INVX1_77/Y OAI22X1_43/D DFFSR_1/gnd NOR2X1_41/B
+ DFFSR_81/S OAI22X1
XFILL_3_NAND3X1_55 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_4_OAI22X1_37 INVX1_3/gnd DFFSR_23/S FILL
XFILL_2_NAND2X1_128 BUFX2_72/gnd DFFSR_276/S FILL
XDFFSR_173 DFFSR_173/Q CLKBUF1_14/Y BUFX2_64/Y DFFSR_208/S DFFSR_165/Q XOR2X1_1/gnd
+ DFFSR_208/S DFFSR
XFILL_2_NAND3X1_58 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_8_DFFSR_32 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_3_OAI22X1_40 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_25_DFFSR_25 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_14_DFFSR_65 BUFX2_79/A DFFSR_7/S FILL
XFILL_4_DFFSR_170 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_1_NAND3X1_61 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_2_OAI22X1_43 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_45_DFFSR_201 INVX1_67/gnd DFFSR_201/S FILL
XFILL_32_6_0 INVX1_1/gnd DFFSR_97/S FILL
XFILL_8_DFFSR_277 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_0_NAND3X1_64 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_21_DFFSR_100 INVX1_1/gnd DFFSR_97/S FILL
XFILL_1_OAI22X1_46 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_35_DFFSR_204 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_0_OAI21X1_110 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_23_DFFPOSX1_40 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_0_AND2X2_14 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_11_DFFSR_103 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_0_OAI22X1_49 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_1_XOR2X1_2 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_25_DFFSR_207 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_49_DFFSR_82 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_7_NAND3X1_243 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_15_DFFSR_210 BUFX2_98/A DFFSR_6/S FILL
XINVX1_66 INVX1_66/A OR2X2_2/gnd INVX1_66/Y DFFSR_216/S INVX1
XFILL_18_CLKBUF1_5 BUFX2_99/A DFFSR_92/S FILL
XFILL_33_DFFSR_32 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_5_DFFSR_79 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_22_DFFSR_72 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_48_DFFSR_128 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_38_DFFSR_131 NOR3X1_6/gnd DFFSR_79/S FILL
XINVX1_184 DFFSR_4/D DFFSR_5/gnd INVX1_184/Y DFFSR_5/S INVX1
XFILL_8_NAND3X1_177 AND2X2_38/B DFFSR_59/S FILL
XCLKBUF1_5 BUFX2_4/Y BUFX2_99/A CLKBUF1_5/Y DFFSR_92/S CLKBUF1
XFILL_1_DFFSR_207 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_4_BUFX2_17 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_28_DFFSR_134 INVX1_1/gnd DFFSR_53/S FILL
XFILL_9_XOR2X1_9 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_42_DFFSR_238 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_1_NAND2X1_158 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_6_NAND3X1_10 BUFX2_79/A DFFSR_6/S FILL
XFILL_4_INVX1_181 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_4_DFFSR_9 BUFX2_79/A DFFSR_6/S FILL
XFILL_4_CLKBUF1_2 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_18_DFFSR_137 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_32_DFFSR_241 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_5_NAND3X1_13 DFFSR_4/gnd DFFSR_4/S FILL
XNAND3X1_10 DFFSR_2/Q NOR2X1_4/Y BUFX2_18/Y BUFX2_79/A AND2X2_7/B DFFSR_6/S NAND3X1
XFILL_22_DFFSR_244 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_4_NAND3X1_16 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_30_DFFSR_79 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_41_DFFSR_39 INVX1_3/gnd DFFSR_79/S FILL
XFILL_2_INVX1_73 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_3_NOR2X1_16 BUFX2_79/A DFFSR_7/S FILL
XFILL_13_DFFPOSX1_15 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_12_DFFSR_247 BUFX2_99/A DFFSR_7/S FILL
XFILL_3_NAND3X1_19 BUFX2_99/A DFFSR_92/S FILL
XDFFSR_137 DFFSR_193/D CLKBUF1_20/Y BUFX2_62/Y DFFSR_216/S INVX1_60/A BUFX2_7/gnd
+ DFFSR_216/S DFFSR
XFILL_42_1_0 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_2_NAND3X1_22 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_14_DFFSR_29 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_4_DFFSR_134 INVX1_1/gnd DFFSR_53/S FILL
XFILL_1_BUFX2_64 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_1_NAND3X1_25 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_45_DFFSR_165 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_8_DFFSR_241 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_0_NAND3X1_28 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_1_OAI22X1_10 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_40_3_1 BUFX2_98/A DFFSR_6/S FILL
XFILL_35_DFFSR_168 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_49_DFFSR_272 INVX1_3/gnd DFFSR_23/S FILL
XFILL_0_OAI22X1_13 INVX1_1/gnd DFFSR_53/S FILL
XFILL_25_DFFSR_171 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_38_DFFSR_86 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_39_DFFSR_275 BUFX2_99/A DFFSR_92/S FILL
XFILL_49_DFFSR_46 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_38_5_2 BUFX2_79/A DFFSR_7/S FILL
XFILL_15_DFFSR_174 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_7_NAND3X1_207 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_7_AOI22X1_6 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_29_DFFSR_278 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_3_DFFPOSX1_26 AND2X2_38/B DFFSR_23/S FILL
XINVX1_30 INVX1_30/A INVX1_1/gnd INVX1_30/Y DFFSR_53/S INVX1
XDFFSR_83 DFFSR_83/Q DFFSR_83/CLK DFFSR_73/R DFFSR_79/S DFFSR_75/Q INVX1_3/gnd DFFSR_79/S
+ DFFSR
XFILL_22_DFFSR_36 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_5_DFFSR_43 BUFX2_98/A DFFSR_6/S FILL
XFILL_11_DFFSR_76 BUFX2_79/A DFFSR_7/S FILL
XFILL_1_XOR2X1_13 INVX1_1/gnd DFFSR_97/S FILL
XFILL_0_NOR2X1_53 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_2_OAI21X1_1 BUFX2_79/A DFFSR_7/S FILL
XINVX1_148 INVX1_148/A BUFX2_7/gnd INVX1_148/Y DFFSR_216/S INVX1
XFILL_8_NAND3X1_141 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_1_DFFSR_171 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_12_DFFPOSX1_45 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_1_NAND2X1_122 INVX1_67/gnd DFFSR_175/S FILL
XFILL_15_XOR2X1_6 BUFX2_99/A DFFSR_7/S FILL
XFILL_42_DFFSR_202 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_49_DFFSR_9 BUFX2_79/A DFFSR_6/S FILL
XFILL_4_INVX1_145 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_46_DFFSR_93 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_7_AND2X2_12 BUFX2_98/A DFFSR_32/S FILL
XFILL_18_DFFSR_101 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_5_DFFSR_278 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_32_DFFSR_205 INVX1_3/gnd DFFSR_79/S FILL
XFILL_7_AND2X2_2 BUFX2_99/A DFFSR_7/S FILL
XFILL_22_DFFSR_208 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_2_DFFSR_90 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_2_INVX1_37 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_30_DFFSR_43 BUFX2_98/A DFFSR_6/S FILL
XFILL_19_DFFSR_83 INVX1_3/gnd DFFSR_79/S FILL
XFILL_12_DFFSR_211 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_22_DFFPOSX1_34 OR2X2_2/gnd DFFSR_216/S FILL
XDFFSR_101 AOI22X1_5/B DFFSR_93/CLK DFFSR_5/R DFFSR_4/S DFFSR_93/Q OR2X2_3/gnd DFFSR_4/S
+ DFFSR
XFILL_15_CLKBUF1_6 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_6_NAND3X1_237 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_1_BUFX2_28 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_45_DFFSR_129 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_8_DFFSR_205 INVX1_3/gnd DFFSR_79/S FILL
XFILL_35_DFFSR_132 INVX1_3/gnd DFFSR_79/S FILL
XFILL_48_0_2 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_49_DFFSR_236 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_25_DFFSR_135 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_49_DFFSR_10 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_1_INVX1_182 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_38_DFFSR_50 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_39_DFFSR_239 INVX1_39/gnd DFFSR_54/S FILL
XFILL_27_DFFSR_90 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_1_CLKBUF1_3 BUFX2_98/A DFFSR_6/S FILL
XFILL_15_DFFSR_138 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_7_NAND3X1_171 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_29_DFFSR_242 OR2X2_3/gnd DFFSR_60/S FILL
XDFFSR_47 DFFSR_63/D CLKBUF1_38/Y DFFSR_15/R DFFSR_98/S DFFSR_39/Q BUFX2_77/gnd DFFSR_98/S
+ DFFSR
XFILL_0_NAND2X1_152 INVX1_1/gnd DFFSR_97/S FILL
XFILL_19_DFFSR_245 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_11_DFFSR_40 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_0_NOR2X1_17 BUFX2_79/A DFFSR_6/S FILL
XFILL_8_NAND3X1_105 DFFSR_1/gnd DFFSR_81/S FILL
XINVX1_112 DFFSR_184/D AND2X2_38/B INVX1_112/Y DFFSR_23/S INVX1
XFILL_1_DFFSR_135 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_15_DFFSR_7 BUFX2_79/A DFFSR_7/S FILL
XFILL_42_DFFSR_166 AND2X2_38/B DFFSR_59/S FILL
XFILL_4_INVX1_109 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_46_DFFSR_57 BUFX2_79/A DFFSR_6/S FILL
XFILL_35_DFFSR_97 INVX1_1/gnd DFFSR_97/S FILL
XFILL_5_DFFSR_242 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_32_DFFSR_169 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_14_1_1 INVX1_39/gnd DFFSR_54/S FILL
XFILL_46_DFFSR_273 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_22_DFFSR_172 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_36_DFFSR_276 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_19_DFFSR_47 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_2_DFFSR_54 INVX1_39/gnd DFFSR_54/S FILL
XFILL_12_DFFSR_175 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_6_BUFX2_82 INVX1_1/gnd DFFSR_97/S FILL
XFILL_4_AOI22X1_7 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_26_DFFSR_279 BUFX2_99/A DFFSR_7/S FILL
XFILL_12_3_2 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_8_XOR2X1_11 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_20_CLKBUF1_37 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_6_NAND3X1_201 INVX1_1/gnd DFFSR_53/S FILL
XFILL_36_DFFSR_3 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_19_CLKBUF1_40 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_2_DFFPOSX1_20 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_8_DFFSR_169 DFFSR_62/gnd DFFSR_62/S FILL
XAND2X2_16 INVX1_62/A NOR3X1_3/A NOR3X1_6/gnd AND2X2_16/Y DFFSR_91/S AND2X2
XFILL_18_CLKBUF1_43 AND2X2_38/B DFFSR_23/S FILL
XFILL_49_DFFSR_200 DFFSR_62/gnd DFFSR_62/S FILL
XNAND3X1_237 XOR2X1_6/Y AOI21X1_37/B AOI21X1_37/A OR2X2_3/gnd NAND3X1_239/A DFFSR_60/S
+ NAND3X1
XFILL_17_CLKBUF1_46 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_38_DFFSR_14 INVX1_1/gnd DFFSR_53/S FILL
XFILL_1_INVX1_146 INVX1_3/gnd DFFSR_79/S FILL
XFILL_39_DFFSR_203 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_4_AND2X2_13 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_16_DFFSR_94 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_27_DFFSR_54 INVX1_39/gnd DFFSR_54/S FILL
XFILL_15_DFFSR_102 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_2_DFFSR_279 BUFX2_99/A DFFSR_7/S FILL
XFILL_7_NAND3X1_135 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_29_DFFSR_206 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_16_CLKBUF1_49 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_11_DFFPOSX1_39 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_19_DFFSR_209 BUFX2_72/gnd DFFSR_276/S FILL
XDFFSR_11 DFFSR_67/D CLKBUF1_8/Y DFFSR_1/R DFFSR_1/S DFFSR_11/D DFFSR_1/gnd DFFSR_1/S
+ DFFSR
XFILL_0_NAND2X1_116 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_39_6_0 BUFX2_79/A DFFSR_6/S FILL
XFILL_12_CLKBUF1_7 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_21_DFFPOSX1_28 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_42_DFFSR_130 BUFX2_79/A DFFSR_6/S FILL
XFILL_35_DFFSR_61 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_46_DFFSR_21 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_5_DFFSR_206 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_32_DFFSR_133 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_46_DFFSR_237 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_5_NAND3X1_231 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_8_CLKBUF1_1 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_22_DFFSR_136 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_1_DFFPOSX1_50 INVX1_1/gnd DFFSR_53/S FILL
XFILL_2_DFFSR_18 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_19_DFFSR_11 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_36_DFFSR_240 INVX1_39/gnd DFFSR_34/S FILL
XFILL_6_BUFX2_46 BUFX2_98/A DFFSR_6/S FILL
XFILL_12_DFFSR_139 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_26_DFFSR_243 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_16_DFFSR_246 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_45_1 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_6_NAND3X1_165 INVX1_39/gnd DFFSR_34/S FILL
XFILL_43_DFFSR_68 BUFX2_98/A DFFSR_6/S FILL
XFILL_8_DFFSR_133 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_49_DFFSR_164 OR2X2_2/gnd DFFSR_216/S FILL
XNAND3X1_201 NAND3X1_201/A OAI21X1_65/Y AOI21X1_30/Y INVX1_1/gnd AOI22X1_26/C DFFSR_53/S
+ NAND3X1
XFILL_17_CLKBUF1_10 INVX1_67/gnd DFFSR_201/S FILL
XFILL_39_DFFSR_167 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_1_INVX1_110 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_16_DFFSR_58 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_27_DFFSR_18 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_2_DFFSR_243 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_3_BUFX2_93 AND2X2_38/B DFFSR_59/S FILL
XFILL_16_CLKBUF1_13 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_29_DFFSR_170 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_43_DFFSR_274 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_15_CLKBUF1_16 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_19_DFFSR_173 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_33_DFFSR_277 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_49_1_0 OR2X2_3/gnd DFFSR_4/S FILL
XNOR2X1_55 NOR2X1_55/A NOR2X1_55/B INVX1_39/gnd NOR2X1_55/Y DFFSR_54/S NOR2X1
XFILL_14_CLKBUF1_19 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_3_DFFSR_6 BUFX2_79/A DFFSR_6/S FILL
XFILL_1_AOI22X1_8 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_23_DFFSR_280 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_51_DFFSR_75 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_5_XOR2X1_12 INVX1_3/gnd DFFSR_23/S FILL
XFILL_13_CLKBUF1_22 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_4_NOR2X1_52 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_47_3_1 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_12_CLKBUF1_25 INVX1_67/gnd DFFSR_201/S FILL
XFILL_7_OAI21X1_117 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_11_CLKBUF1_28 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_7_DFFSR_72 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_35_DFFSR_25 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_24_DFFSR_65 BUFX2_79/A DFFSR_7/S FILL
XFILL_5_DFFSR_170 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_10_CLKBUF1_31 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_46_DFFSR_201 INVX1_67/gnd DFFSR_201/S FILL
XFILL_45_5_2 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_5_NAND3X1_195 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_9_DFFSR_277 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_22_DFFSR_100 INVX1_1/gnd DFFSR_97/S FILL
XFILL_36_DFFSR_204 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_1_OR2X2_6 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_1_DFFPOSX1_14 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_1_AND2X2_14 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_12_DFFSR_103 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_9_CLKBUF1_34 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_26_DFFSR_207 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_16_DFFSR_210 BUFX2_98/A DFFSR_6/S FILL
XFILL_8_CLKBUF1_37 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_6_NAND3X1_129 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_7_CLKBUF1_40 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_19_CLKBUF1_5 BUFX2_99/A DFFSR_92/S FILL
XFILL_10_DFFPOSX1_33 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_4_INVX1_66 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_43_DFFSR_32 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_32_DFFSR_72 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_6_CLKBUF1_43 AND2X2_38/B DFFSR_23/S FILL
XFILL_49_DFFSR_128 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_13_4_0 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_5_CLKBUF1_46 OR2X2_3/gnd DFFSR_4/S FILL
XNAND3X1_165 AOI21X1_13/A OAI21X1_41/Y AOI21X1_13/C INVX1_39/gnd AOI21X1_26/C DFFSR_34/S
+ NAND3X1
XFILL_39_DFFSR_131 NOR3X1_6/gnd DFFSR_79/S FILL
XCLKBUF1_43 clk AND2X2_38/B CLKBUF1_43/Y DFFSR_23/S CLKBUF1
XFILL_16_DFFSR_22 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_4_CLKBUF1_49 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_2_DFFSR_207 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_3_BUFX2_57 AND2X2_38/B DFFSR_23/S FILL
XFILL_29_DFFSR_134 INVX1_1/gnd DFFSR_53/S FILL
XFILL_11_6_1 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_43_DFFSR_238 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_20_DFFPOSX1_22 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_5_CLKBUF1_2 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_19_DFFSR_137 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_33_DFFSR_241 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_7_NOR3X1_3 BUFX2_7/gnd DFFSR_216/S FILL
XNOR2X1_19 NOR2X1_19/A NOR2X1_19/B DFFSR_28/gnd NOR2X1_19/Y DFFSR_3/S NOR2X1
XFILL_48_DFFSR_6 BUFX2_79/A DFFSR_6/S FILL
XFILL_23_DFFSR_244 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_4_NAND3X1_225 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_40_DFFSR_79 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_51_DFFSR_39 INVX1_3/gnd DFFSR_79/S FILL
XFILL_4_NOR2X1_16 BUFX2_79/A DFFSR_7/S FILL
XFILL_13_DFFSR_247 BUFX2_99/A DFFSR_7/S FILL
XFILL_0_DFFPOSX1_44 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_50_6 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_24_DFFSR_29 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_7_DFFSR_36 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_13_DFFSR_69 BUFX2_98/A DFFSR_32/S FILL
XFILL_5_DFFSR_134 INVX1_1/gnd DFFSR_53/S FILL
XFILL_46_DFFSR_165 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_5_NAND3X1_159 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_9_DFFSR_241 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_36_DFFSR_168 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_3_INVX1_8 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_50_DFFSR_272 INVX1_3/gnd DFFSR_23/S FILL
XFILL_0_XOR2X1_6 BUFX2_99/A DFFSR_7/S FILL
XFILL_26_DFFSR_171 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_40_DFFSR_275 BUFX2_99/A DFFSR_92/S FILL
XFILL_48_DFFSR_86 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_16_DFFSR_174 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_8_AOI22X1_6 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_30_DFFSR_278 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_4_DFFSR_83 INVX1_3/gnd DFFSR_79/S FILL
XFILL_32_DFFSR_36 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_21_DFFSR_76 BUFX2_79/A DFFSR_7/S FILL
XFILL_2_XOR2X1_13 INVX1_1/gnd DFFSR_97/S FILL
XFILL_1_NOR2X1_53 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_3_OAI21X1_1 BUFX2_79/A DFFSR_7/S FILL
XFILL_5_CLKBUF1_10 INVX1_67/gnd DFFSR_201/S FILL
XNAND3X1_129 AOI21X1_1/A AOI21X1_1/B INVX1_120/A DFFSR_62/gnd AND2X2_27/B DFFSR_62/S
+ NAND3X1
XFILL_21_1_1 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_4_CLKBUF1_13 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_2_DFFSR_171 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_3_BUFX2_21 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_3_0_0 INVX1_67/gnd DFFSR_175/S FILL
XFILL_3_CLKBUF1_16 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_43_DFFSR_202 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_8_AND2X2_12 BUFX2_98/A DFFSR_32/S FILL
XFILL_19_DFFSR_101 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_6_OAI21X1_111 AND2X2_38/B DFFSR_59/S FILL
XFILL_19_3_2 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_6_DFFSR_278 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_33_DFFSR_205 INVX1_3/gnd DFFSR_79/S FILL
XFILL_2_CLKBUF1_19 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_14_DFFSR_4 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_1_2_1 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_4_NAND3X1_189 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_23_DFFSR_208 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_1_CLKBUF1_22 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_40_DFFSR_43 BUFX2_98/A DFFSR_6/S FILL
XFILL_29_DFFSR_83 INVX1_3/gnd DFFSR_79/S FILL
XFILL_1_INVX1_77 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_13_DFFSR_211 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_0_CLKBUF1_25 INVX1_67/gnd DFFSR_201/S FILL
XFILL_16_CLKBUF1_6 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_13_DFFSR_33 BUFX2_98/A DFFSR_32/S FILL
XFILL_0_BUFX2_68 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_46_DFFSR_129 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_5_NAND3X1_123 BUFX2_99/A DFFSR_7/S FILL
XFILL_9_DFFSR_205 INVX1_3/gnd DFFSR_79/S FILL
XFILL_36_DFFSR_132 INVX1_3/gnd DFFSR_79/S FILL
XFILL_50_DFFSR_236 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_26_DFFSR_135 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_10_3 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_2_INVX1_182 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_48_DFFSR_50 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_40_DFFSR_239 INVX1_39/gnd DFFSR_54/S FILL
XFILL_37_DFFSR_90 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_2_CLKBUF1_3 BUFX2_98/A DFFSR_6/S FILL
XFILL_16_DFFSR_138 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_46_6_0 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_30_DFFSR_242 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_20_DFFSR_245 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_4_DFFSR_47 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_19_DFFPOSX1_16 INVX1_67/gnd DFFSR_175/S FILL
XFILL_21_DFFSR_40 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_10_DFFSR_80 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_1_NOR2X1_17 BUFX2_79/A DFFSR_6/S FILL
XFILL_10_DFFSR_248 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_3_NAND3X1_219 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_2_DFFSR_135 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_27_DFFPOSX1_4 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_43_DFFSR_166 AND2X2_38/B DFFSR_59/S FILL
XFILL_45_DFFSR_97 INVX1_1/gnd DFFSR_97/S FILL
XFILL_6_DFFSR_242 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_26_DFFPOSX1_7 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_33_DFFSR_169 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_47_DFFSR_273 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_6_AND2X2_6 BUFX2_99/A DFFSR_7/S FILL
XFILL_23_DFFSR_172 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_4_NAND3X1_153 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_37_DFFSR_276 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_1_INVX1_41 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_29_DFFSR_47 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_1_DFFSR_94 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_18_DFFSR_87 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_13_DFFSR_175 OR2X2_2/gnd DFFSR_175/S FILL
XOAI21X1_111 NAND3X1_8/Y NAND3X1_72/Y INVX1_212/Y AND2X2_38/B NOR2X1_77/B DFFSR_59/S
+ OAI21X1
XFILL_5_AOI22X1_7 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_27_DFFSR_279 BUFX2_99/A DFFSR_7/S FILL
XFILL_9_DFFPOSX1_27 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_9_XOR2X1_11 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_0_BUFX2_32 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_0_OAI21X1_2 BUFX2_79/A DFFSR_7/S FILL
XFILL_9_DFFSR_169 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_18_DFFPOSX1_46 INVX1_39/gnd DFFSR_34/S FILL
XFILL_50_DFFSR_200 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_48_DFFSR_14 INVX1_1/gnd DFFSR_53/S FILL
XFILL_2_INVX1_146 INVX1_3/gnd DFFSR_79/S FILL
XFILL_40_DFFSR_203 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_5_AND2X2_13 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_26_DFFSR_94 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_37_DFFSR_54 INVX1_39/gnd DFFSR_54/S FILL
XFILL_16_DFFSR_102 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_2_NAND3X1_249 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_3_DFFSR_279 BUFX2_99/A DFFSR_7/S FILL
XFILL_30_DFFSR_206 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_54_3_1 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_20_DFFSR_209 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_4_DFFSR_11 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_10_DFFSR_44 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_5_OAI21X1_105 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_10_DFFSR_212 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_52_5_2 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_3_NAND3X1_183 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_13_CLKBUF1_7 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_2_DFFSR_3 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_43_DFFSR_130 BUFX2_79/A DFFSR_6/S FILL
XFILL_45_DFFSR_61 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_6_DFFSR_206 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_33_DFFSR_133 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_47_DFFSR_237 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_9_CLKBUF1_1 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_23_DFFSR_136 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_4_NAND3X1_117 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_1_DFFSR_58 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_29_DFFSR_11 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_37_DFFSR_240 INVX1_39/gnd DFFSR_34/S FILL
XFILL_18_DFFSR_51 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_13_DFFSR_139 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_5_BUFX2_86 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_27_DFFSR_243 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_6_NAND2X1_153 BUFX2_98/A DFFSR_32/S FILL
XFILL_32_3 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_0_OR2X2_3 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_20_4_0 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_17_DFFSR_246 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_9_DFFSR_133 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_26_DFFSR_7 BUFX2_79/A DFFSR_7/S FILL
XFILL_18_6_1 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_18_DFFPOSX1_10 INVX1_67/gnd DFFSR_201/S FILL
XFILL_50_DFFSR_164 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_0_5_0 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_40_DFFSR_167 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_9_DFFSR_65 BUFX2_79/A DFFSR_7/S FILL
XFILL_2_INVX1_110 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_26_DFFSR_58 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_15_DFFSR_98 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_37_DFFSR_18 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_2_NAND3X1_213 INVX1_39/gnd DFFSR_54/S FILL
XFILL_3_DFFSR_243 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_30_DFFSR_170 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_44_DFFSR_274 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_20_DFFSR_173 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_34_DFFSR_277 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_16_DFFPOSX1_1 INVX1_39/gnd DFFSR_34/S FILL
XFILL_10_DFFSR_176 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_2_AOI22X1_8 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_24_DFFSR_280 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_15_DFFPOSX1_4 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_6_XOR2X1_12 INVX1_3/gnd DFFSR_23/S FILL
XFILL_3_NAND3X1_147 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_5_NOR2X1_52 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_47_DFFSR_3 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_14_DFFPOSX1_7 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_8_DFFPOSX1_21 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_45_DFFSR_25 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_34_DFFSR_65 BUFX2_79/A DFFSR_7/S FILL
XFILL_6_DFFSR_170 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_47_DFFSR_201 INVX1_67/gnd DFFSR_201/S FILL
XFILL_23_DFFSR_100 INVX1_1/gnd DFFSR_97/S FILL
XFILL_37_DFFSR_204 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_1_DFFSR_22 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_18_DFFSR_15 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_2_AND2X2_14 DFFSR_46/gnd DFFSR_54/S FILL
XBUFX2_90 BUFX2_90/A OR2X2_2/gnd BUFX2_90/Y DFFSR_175/S BUFX2
XFILL_13_DFFSR_103 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_5_BUFX2_50 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_0_DFFSR_280 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_17_DFFPOSX1_40 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_27_DFFSR_207 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_6_NAND2X1_117 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_2_INVX1_5 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_17_DFFSR_210 BUFX2_98/A DFFSR_6/S FILL
XFILL_28_1_1 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_1_NAND3X1_243 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_0_NOR2X1_3 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_20_CLKBUF1_5 BUFX2_99/A DFFSR_92/S FILL
XFILL_42_DFFSR_72 OR2X2_3/gnd DFFSR_60/S FILL
XNAND2X1_153 DFFSR_6/S NAND2X1_153/B BUFX2_98/A AOI21X1_52/B DFFSR_32/S NAND2X1
XFILL_10_CLKBUF1_8 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_50_DFFSR_128 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_26_3_2 INVX1_3/gnd DFFSR_23/S FILL
XFILL_27_DFFPOSX1_29 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_8_AOI21X1_45 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_8_2_1 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_9_DFFSR_29 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_40_DFFSR_131 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_26_DFFSR_22 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_7_AOI21X1_48 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_15_DFFSR_62 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_2_NAND3X1_177 AND2X2_38/B DFFSR_59/S FILL
XFILL_3_DFFSR_207 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_2_BUFX2_97 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_30_DFFSR_134 INVX1_1/gnd DFFSR_53/S FILL
XFILL_6_AOI21X1_51 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_44_DFFSR_238 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_6_CLKBUF1_2 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_20_DFFSR_137 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_6_4_2 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_5_AOI21X1_54 AND2X2_38/B DFFSR_59/S FILL
XFILL_34_DFFSR_241 BUFX2_72/gnd DFFSR_201/S FILL
XAOI21X1_51 AOI21X1_51/A AOI21X1_51/B BUFX2_35/Y DFFSR_1/gnd AOI21X1_51/Y DFFSR_81/S
+ AOI21X1
XFILL_10_DFFSR_140 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_4_AOI21X1_57 INVX1_67/gnd DFFSR_201/S FILL
XFILL_24_DFFSR_244 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_50_DFFSR_79 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_3_NAND3X1_111 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_5_NOR2X1_16 BUFX2_79/A DFFSR_7/S FILL
XFILL_13_DFFSR_1 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_3_AOI21X1_60 BUFX2_79/A DFFSR_7/S FILL
XFILL_14_DFFSR_247 BUFX2_99/A DFFSR_7/S FILL
XFILL_2_AOI21X1_63 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_54_3 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_5_NAND2X1_147 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_34_DFFSR_29 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_6_DFFSR_76 BUFX2_79/A DFFSR_7/S FILL
XFILL_23_DFFSR_69 BUFX2_98/A DFFSR_32/S FILL
XFILL_6_DFFSR_134 INVX1_1/gnd DFFSR_53/S FILL
XFILL_1_AOI21X1_66 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_47_DFFSR_165 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_53_6_0 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_0_AOI21X1_69 INVX1_1/gnd DFFSR_97/S FILL
XFILL_37_DFFSR_168 OR2X2_6/gnd DFFSR_92/S FILL
XBUFX2_54 BUFX2_53/A BUFX2_7/gnd BUFX2_54/Y DFFSR_151/S BUFX2
XFILL_5_BUFX2_14 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_0_DFFSR_244 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_27_DFFSR_171 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_41_DFFSR_275 BUFX2_99/A DFFSR_92/S FILL
XFILL_17_DFFSR_174 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_8_OAI21X1_93 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_9_AOI22X1_6 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_31_DFFSR_278 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_1_NAND3X1_207 DFFSR_1/gnd DFFSR_1/S FILL
XOAI21X1_4 INVX1_30/Y OAI21X1_4/B OAI21X1_4/C OR2X2_6/gnd OAI21X1_4/Y DFFSR_53/S OAI21X1
XFILL_7_OAI21X1_96 AND2X2_38/B DFFSR_59/S FILL
XFILL_42_DFFSR_36 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_31_DFFSR_76 BUFX2_79/A DFFSR_7/S FILL
XFILL_3_INVX1_70 NOR3X1_6/gnd DFFSR_79/S FILL
XNAND2X1_117 DFFSR_98/S din[1] BUFX2_77/gnd OAI21X1_86/C DFFSR_5/S NAND2X1
XFILL_3_XOR2X1_13 INVX1_1/gnd DFFSR_97/S FILL
XFILL_2_NOR2X1_53 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_6_OAI21X1_99 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_4_OAI21X1_1 BUFX2_79/A DFFSR_7/S FILL
XFILL_15_DFFSR_26 BUFX2_79/A DFFSR_6/S FILL
XFILL_7_AOI21X1_12 DFFSR_1/gnd DFFSR_1/S FILL
XOAI21X1_99 BUFX2_52/Y INVX1_196/Y OAI21X1_99/C DFFSR_34/gnd DFFSR_271/D DFFSR_1/S
+ OAI21X1
XFILL_3_DFFSR_171 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_2_NAND3X1_141 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_2_BUFX2_61 AND2X2_38/B DFFSR_59/S FILL
XFILL_6_AOI21X1_15 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_44_DFFSR_202 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_7_DFFPOSX1_15 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_20_DFFSR_101 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_5_AOI21X1_18 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_4_DFFPOSX1_1 INVX1_39/gnd DFFSR_34/S FILL
XFILL_7_DFFSR_278 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_4_NAND2X1_177 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_34_DFFSR_205 INVX1_3/gnd DFFSR_79/S FILL
XFILL_10_DFFSR_104 DFFSR_28/gnd DFFSR_8/S FILL
XAOI21X1_15 INVX1_143/Y AOI21X1_15/B AOI21X1_15/C DFFSR_1/gnd AOI21X1_15/Y DFFSR_81/S
+ AOI21X1
XFILL_3_DFFPOSX1_4 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_4_AOI21X1_21 INVX1_39/gnd DFFSR_54/S FILL
XFILL_24_DFFSR_208 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_50_DFFSR_43 BUFX2_98/A DFFSR_6/S FILL
XFILL_39_DFFSR_83 INVX1_3/gnd DFFSR_79/S FILL
XFILL_2_DFFPOSX1_7 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_3_AOI21X1_24 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_14_DFFSR_211 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_16_DFFPOSX1_34 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_2_AOI21X1_27 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_17_CLKBUF1_6 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_6_DFFSR_40 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_5_NAND2X1_111 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_23_DFFSR_33 BUFX2_98/A DFFSR_32/S FILL
XFILL_1_AOI21X1_30 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_12_DFFSR_73 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_47_DFFSR_129 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_0_NAND3X1_237 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_0_AOI21X1_33 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_37_DFFSR_132 INVX1_3/gnd DFFSR_79/S FILL
XBUFX2_18 NOR2X1_7/Y BUFX2_98/A BUFX2_18/Y DFFSR_32/S BUFX2
XFILL_0_DFFSR_208 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_27_DFFSR_135 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_16_XOR2X1_3 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_9_OAI21X1_54 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_3_INVX1_182 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_26_DFFPOSX1_23 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_41_DFFSR_239 INVX1_39/gnd DFFSR_54/S FILL
XFILL_47_DFFSR_90 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_3_CLKBUF1_3 BUFX2_98/A DFFSR_6/S FILL
XFILL_17_DFFSR_138 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_31_DFFSR_242 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_8_OAI21X1_57 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_1_NAND3X1_171 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_6_NAND2X1_78 AND2X2_38/B DFFSR_23/S FILL
XFILL_7_OAI21X1_60 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_21_DFFSR_245 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_31_DFFSR_40 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_20_DFFSR_80 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_3_DFFSR_87 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_3_INVX1_34 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_2_NOR2X1_17 BUFX2_79/A DFFSR_6/S FILL
XFILL_6_DFFPOSX1_45 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_6_OAI21X1_63 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_5_NAND2X1_81 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_11_DFFSR_248 DFFSR_28/gnd DFFSR_8/S FILL
XNAND2X1_78 NAND2X1_77/B AND2X2_34/Y AND2X2_38/B NAND2X1_78/Y DFFSR_23/S NAND2X1
XFILL_5_OAI21X1_66 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_4_NAND2X1_84 NOR3X1_6/gnd DFFSR_91/S FILL
XOAI21X1_63 XNOR2X1_3/A INVX1_166/Y OAI21X1_62/Y XOR2X1_4/gnd OAI21X1_63/Y DFFSR_97/S
+ OAI21X1
XFILL_2_NAND3X1_105 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_3_DFFSR_135 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_3_NAND2X1_87 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_4_OAI21X1_69 INVX1_3/gnd DFFSR_23/S FILL
XFILL_2_BUFX2_25 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_44_DFFSR_166 AND2X2_38/B DFFSR_59/S FILL
XFILL_3_OAI21X1_72 INVX1_3/gnd DFFSR_23/S FILL
XFILL_2_NAND2X1_90 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_7_DFFSR_242 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_27_4_0 INVX1_3/gnd DFFSR_79/S FILL
XFILL_4_NAND2X1_141 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_34_DFFSR_169 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_1_NAND2X1_93 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_12_NOR3X1_4 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_2_OAI21X1_75 INVX1_39/gnd DFFSR_54/S FILL
XFILL_48_DFFSR_273 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_24_DFFSR_172 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_0_NAND2X1_96 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_38_DFFSR_276 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_1_OAI21X1_78 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_0_INVX1_81 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_28_DFFSR_87 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_39_DFFSR_47 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_14_DFFSR_175 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_25_6_1 AND2X2_38/B DFFSR_23/S FILL
XFILL_6_AOI22X1_7 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_0_OAI21X1_81 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_28_DFFSR_279 BUFX2_99/A DFFSR_7/S FILL
XFILL_7_5_0 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_12_DFFSR_37 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_0_XOR2X1_14 INVX1_1/gnd DFFSR_53/S FILL
XFILL_0_NAND3X1_201 INVX1_1/gnd DFFSR_53/S FILL
XFILL_1_OAI21X1_2 BUFX2_79/A DFFSR_7/S FILL
XFILL_0_DFFSR_172 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_25_DFFSR_4 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_3_INVX1_146 INVX1_3/gnd DFFSR_79/S FILL
XFILL_41_DFFSR_203 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_6_AND2X2_13 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_36_DFFSR_94 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_47_DFFSR_54 INVX1_39/gnd DFFSR_54/S FILL
XFILL_17_DFFSR_102 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_4_DFFSR_279 BUFX2_99/A DFFSR_7/S FILL
XFILL_31_DFFSR_206 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_8_OAI21X1_21 AND2X2_38/B DFFSR_59/S FILL
XFILL_1_NAND3X1_135 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_21_DFFSR_209 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_7_OAI21X1_24 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_6_NAND2X1_42 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_20_DFFSR_44 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_3_DFFSR_51 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_6_OAI21X1_27 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_3_NAND2X1_171 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_5_NAND2X1_45 INVX1_39/gnd DFFSR_34/S FILL
XFILL_11_DFFSR_212 OR2X2_2/gnd DFFSR_175/S FILL
XNAND2X1_42 DFFSR_163/Q AND2X2_18/Y DFFSR_34/gnd NAND3X1_84/A DFFSR_34/S NAND2X1
XFILL_4_NAND2X1_48 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_5_OAI21X1_30 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_14_CLKBUF1_7 OR2X2_4/gnd DFFSR_32/S FILL
XOAI21X1_27 NOR2X1_68/Y AND2X2_30/Y INVX1_131/Y OR2X2_2/gnd OAI21X1_27/Y DFFSR_216/S
+ OAI21X1
XFILL_3_NAND2X1_51 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_4_OAI21X1_33 INVX1_3/gnd DFFSR_79/S FILL
XDFFPOSX1_45 INVX1_145/A CLKBUF1_48/Y AOI21X1_64/Y OR2X2_1/gnd DFFSR_59/S DFFPOSX1
XFILL_44_DFFSR_130 BUFX2_79/A DFFSR_6/S FILL
XFILL_15_DFFPOSX1_28 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_2_NAND2X1_54 AND2X2_38/B DFFSR_59/S FILL
XFILL_3_OAI21X1_36 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_7_DFFSR_206 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_34_DFFSR_133 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_4_NAND2X1_105 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_1_NAND2X1_57 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_2_OAI21X1_39 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_48_DFFSR_237 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_35_1_1 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_24_DFFSR_136 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_0_NAND2X1_60 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_1_OAI21X1_42 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_0_INVX1_45 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_0_INVX1_183 BUFX2_79/A DFFSR_6/S FILL
XFILL_39_DFFSR_11 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_38_DFFSR_240 INVX1_39/gnd DFFSR_34/S FILL
XFILL_0_DFFSR_98 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_17_DFFSR_91 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_28_DFFSR_51 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_0_CLKBUF1_4 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_14_DFFSR_139 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_19_5 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_28_DFFSR_243 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_0_OAI21X1_45 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_33_3_2 INVX1_1/gnd DFFSR_53/S FILL
XFILL_9_AOI22X1_11 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_25_DFFPOSX1_17 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_18_DFFSR_246 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_0_NAND3X1_165 INVX1_39/gnd DFFSR_34/S FILL
XFILL_8_AOI22X1_14 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_1_INVX1_2 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_9_NAND3X1_220 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_7_AOI22X1_17 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_51_DFFSR_164 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_5_DFFPOSX1_39 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_0_DFFSR_136 NOR3X1_6/gnd DFFSR_79/S FILL
XDFFSR_246 DFFSR_246/Q CLKBUF1_11/Y BUFX2_67/Y DFFSR_208/S DFFSR_238/Q XOR2X1_1/gnd
+ DFFSR_208/S DFFSR
XFILL_6_AOI22X1_20 INVX1_39/gnd DFFSR_34/S FILL
XFILL_41_DFFSR_167 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_3_INVX1_110 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_36_DFFSR_58 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_47_DFFSR_18 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_25_DFFSR_98 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_5_AOI22X1_23 INVX1_39/gnd DFFSR_34/S FILL
XFILL_4_DFFSR_243 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_31_DFFSR_170 OR2X2_6/gnd DFFSR_92/S FILL
XAOI22X1_20 AOI22X1_20/A AOI21X1_9/A AOI22X1_20/C AOI22X1_20/D INVX1_39/gnd NOR3X1_5/B
+ DFFSR_34/S AOI22X1
XFILL_45_DFFSR_274 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_4_AOI22X1_26 INVX1_1/gnd DFFSR_97/S FILL
XFILL_21_DFFSR_173 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_35_DFFSR_277 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_3_DFFSR_15 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_3_AOI22X1_29 INVX1_1/gnd DFFSR_53/S FILL
XFILL_3_NAND2X1_135 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_11_DFFSR_176 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_3_AOI22X1_8 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_25_DFFSR_280 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_4_NAND2X1_12 INVX1_3/gnd DFFSR_79/S FILL
XFILL_7_XOR2X1_12 INVX1_3/gnd DFFSR_23/S FILL
XFILL_6_NOR2X1_52 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_3_NAND2X1_15 BUFX2_99/A DFFSR_92/S FILL
XFILL_2_NAND2X1_18 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_44_DFFSR_65 BUFX2_79/A DFFSR_7/S FILL
XFILL_7_DFFSR_170 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_1_OAI21X1_117 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_24_DFFPOSX1_47 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_1_NAND2X1_21 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_48_DFFSR_201 INVX1_67/gnd DFFSR_201/S FILL
XFILL_8_NAND3X1_77 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_24_DFFSR_100 INVX1_1/gnd DFFSR_97/S FILL
XFILL_0_NAND2X1_24 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_38_DFFSR_204 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_0_INVX1_147 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_0_DFFSR_62 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_28_DFFSR_15 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_17_DFFSR_55 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_3_AND2X2_14 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_14_DFFSR_103 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_4_BUFX2_90 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_1_DFFSR_280 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_7_NAND3X1_80 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_28_DFFSR_207 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_6_NAND3X1_83 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_18_DFFSR_210 BUFX2_98/A DFFSR_6/S FILL
XFILL_5_NAND3X1_86 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_0_NAND3X1_129 DFFSR_62/gnd DFFSR_62/S FILL
XNAND3X1_83 BUFX2_92/A AND2X2_16/Y BUFX2_31/Y XOR2X1_1/gnd AND2X2_21/A DFFSR_151/S
+ NAND3X1
XFILL_4_NAND3X1_89 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_11_CLKBUF1_8 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_0_DFFSR_100 INVX1_1/gnd DFFSR_97/S FILL
XFILL_3_NAND3X1_92 DFFSR_34/gnd DFFSR_1/S FILL
XDFFSR_210 INVX1_71/A DFFSR_3/CLK BUFX2_65/Y DFFSR_6/S INVX1_72/A BUFX2_98/A DFFSR_6/S
+ DFFSR
XFILL_2_NAND2X1_165 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_41_DFFSR_131 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_2_NAND3X1_95 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_36_DFFSR_22 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_8_DFFSR_69 BUFX2_98/A DFFSR_32/S FILL
XFILL_25_DFFSR_62 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_4_DFFSR_207 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_31_DFFSR_134 INVX1_1/gnd DFFSR_53/S FILL
XFILL_1_NAND3X1_98 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_45_DFFSR_238 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_7_CLKBUF1_2 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_21_DFFSR_137 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_35_DFFSR_241 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_14_DFFPOSX1_22 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_11_DFFSR_140 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_25_DFFSR_244 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_6_NOR2X1_16 BUFX2_79/A DFFSR_7/S FILL
XFILL_11_OAI22X1_17 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_37_DFFSR_7 BUFX2_79/A DFFSR_7/S FILL
XFILL_15_DFFSR_247 BUFX2_99/A DFFSR_7/S FILL
XFILL_10_OAI22X1_20 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_44_DFFSR_29 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_33_DFFSR_69 BUFX2_98/A DFFSR_32/S FILL
XFILL_7_DFFSR_134 INVX1_1/gnd DFFSR_53/S FILL
XFILL_24_DFFPOSX1_11 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_9_NAND3X1_38 BUFX2_98/A DFFSR_32/S FILL
XFILL_48_DFFSR_165 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_8_NAND3X1_41 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_9_OAI22X1_23 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_0_DFFSR_26 BUFX2_79/A DFFSR_6/S FILL
XFILL_38_DFFSR_168 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_0_INVX1_111 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_8_NAND3X1_214 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_17_DFFSR_19 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_4_BUFX2_54 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_7_NAND3X1_44 BUFX2_99/A DFFSR_7/S FILL
XFILL_1_DFFSR_244 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_8_OAI22X1_26 INVX1_39/gnd DFFSR_54/S FILL
XFILL_4_DFFPOSX1_33 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_28_DFFSR_171 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_42_DFFSR_275 BUFX2_99/A DFFSR_92/S FILL
XFILL_6_NAND3X1_47 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_7_OAI22X1_29 INVX1_3/gnd DFFSR_79/S FILL
XFILL_18_DFFSR_174 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_32_DFFSR_278 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_5_NAND3X1_50 BUFX2_98/A DFFSR_6/S FILL
XFILL_6_OAI22X1_32 INVX1_39/gnd DFFSR_54/S FILL
XNAND3X1_47 NAND3X1_45/Y NAND3X1_47/B AOI22X1_6/Y OR2X2_3/gnd NOR2X1_23/B DFFSR_4/S
+ NAND3X1
XFILL_0_AOI22X1_9 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_9_NAND3X1_148 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_4_NAND3X1_53 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_41_DFFSR_76 BUFX2_79/A DFFSR_7/S FILL
XFILL_5_OAI22X1_35 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_4_XOR2X1_13 INVX1_1/gnd DFFSR_97/S FILL
XFILL_3_NOR2X1_53 DFFSR_1/gnd DFFSR_81/S FILL
XOAI22X1_32 INVX1_78/Y OAI22X1_41/B INVX1_79/Y OAI22X1_41/D INVX1_39/gnd NOR2X1_41/A
+ DFFSR_54/S OAI22X1
XFILL_3_NAND3X1_56 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_5_OAI21X1_1 BUFX2_79/A DFFSR_7/S FILL
XFILL_4_OAI22X1_38 AND2X2_38/B DFFSR_23/S FILL
XFILL_34_4_0 OR2X2_6/gnd DFFSR_53/S FILL
XDFFSR_174 DFFSR_190/D CLKBUF1_17/Y BUFX2_61/Y DFFSR_51/S DFFSR_174/D BUFX2_8/gnd
+ DFFSR_51/S DFFSR
XFILL_2_NAND2X1_129 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_2_NAND3X1_59 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_3_OAI22X1_41 INVX1_39/gnd DFFSR_54/S FILL
XFILL_8_DFFSR_33 BUFX2_98/A DFFSR_32/S FILL
XFILL_25_DFFSR_26 BUFX2_79/A DFFSR_6/S FILL
XFILL_14_DFFSR_66 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_4_DFFSR_171 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_1_NAND3X1_62 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_2_OAI22X1_44 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_32_6_1 INVX1_1/gnd DFFSR_97/S FILL
XFILL_45_DFFSR_202 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_21_DFFSR_101 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_1_OAI22X1_47 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_0_NAND3X1_65 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_8_DFFSR_278 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_35_DFFSR_205 INVX1_3/gnd DFFSR_79/S FILL
XFILL_0_OAI21X1_111 AND2X2_38/B DFFSR_59/S FILL
XFILL_23_DFFPOSX1_41 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_0_AND2X2_15 INVX1_3/gnd DFFSR_23/S FILL
XFILL_11_DFFSR_104 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_0_OAI22X1_50 INVX1_3/gnd DFFSR_23/S FILL
XFILL_1_XOR2X1_3 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_25_DFFSR_208 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_49_DFFSR_83 INVX1_3/gnd DFFSR_79/S FILL
XFILL_15_DFFSR_211 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_7_NAND3X1_244 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_18_CLKBUF1_6 OR2X2_1/gnd DFFSR_51/S FILL
XINVX1_67 INVX1_67/A INVX1_67/gnd INVX1_67/Y DFFSR_201/S INVX1
XFILL_5_DFFSR_80 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_33_DFFSR_33 BUFX2_98/A DFFSR_32/S FILL
XFILL_22_DFFSR_73 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_48_DFFSR_129 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_8_NAND3X1_178 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_38_DFFSR_132 INVX1_3/gnd DFFSR_79/S FILL
XINVX1_185 DFFSR_5/D DFFSR_4/gnd INVX1_185/Y DFFSR_4/S INVX1
XCLKBUF1_6 BUFX2_5/Y OR2X2_1/gnd CLKBUF1_6/Y DFFSR_51/S CLKBUF1
XFILL_4_BUFX2_18 BUFX2_98/A DFFSR_32/S FILL
XFILL_1_DFFSR_208 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_28_DFFSR_135 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_4_INVX1_182 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_1_NAND2X1_159 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_42_DFFSR_239 INVX1_39/gnd DFFSR_54/S FILL
XFILL_6_NAND3X1_11 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_4_CLKBUF1_3 BUFX2_98/A DFFSR_6/S FILL
XFILL_18_DFFSR_138 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_32_DFFSR_242 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_5_NAND3X1_14 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_24_DFFSR_1 DFFSR_1/gnd DFFSR_1/S FILL
XNAND3X1_11 BUFX2_83/A AND2X2_3/Y BUFX2_21/Y OR2X2_4/gnd AND2X2_7/A DFFSR_32/S NAND3X1
XFILL_4_NAND3X1_17 BUFX2_99/A DFFSR_7/S FILL
XFILL_9_NAND3X1_112 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_22_DFFSR_245 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_41_DFFSR_40 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_2_INVX1_74 BUFX2_99/A DFFSR_92/S FILL
XFILL_30_DFFSR_80 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_3_NOR2X1_17 BUFX2_79/A DFFSR_6/S FILL
XFILL_13_DFFPOSX1_16 INVX1_67/gnd DFFSR_175/S FILL
XFILL_12_DFFSR_248 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_3_NAND3X1_20 BUFX2_99/A DFFSR_7/S FILL
XDFFSR_138 DFFSR_194/D CLKBUF1_6/Y BUFX2_70/Y DFFSR_81/S INVX1_69/A BUFX2_8/gnd DFFSR_81/S
+ DFFSR
XFILL_42_1_1 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_2_NAND3X1_23 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_14_DFFSR_30 BUFX2_98/A DFFSR_32/S FILL
XFILL_4_DFFSR_135 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_1_NAND3X1_26 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_1_BUFX2_65 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_45_DFFSR_166 AND2X2_38/B DFFSR_59/S FILL
XFILL_8_DFFSR_242 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_0_NAND3X1_29 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_40_3_2 BUFX2_98/A DFFSR_6/S FILL
XFILL_1_OAI22X1_11 BUFX2_99/A DFFSR_92/S FILL
XFILL_35_DFFSR_169 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_49_DFFSR_273 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_0_OAI22X1_14 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_25_DFFSR_172 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_39_DFFSR_276 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_38_DFFSR_87 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_49_DFFSR_47 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_15_DFFSR_175 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_7_NAND3X1_208 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_7_AOI22X1_7 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_29_DFFSR_279 BUFX2_99/A DFFSR_7/S FILL
XFILL_3_DFFPOSX1_27 DFFSR_34/gnd DFFSR_1/S FILL
XDFFSR_84 INVX1_26/A DFFSR_92/CLK DFFSR_7/R DFFSR_7/S DFFSR_84/D BUFX2_99/A DFFSR_7/S
+ DFFSR
XINVX1_31 INVX1_31/A INVX1_1/gnd INVX1_31/Y DFFSR_53/S INVX1
XFILL_22_DFFSR_37 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_5_DFFSR_44 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_11_DFFSR_77 BUFX2_98/A DFFSR_32/S FILL
XFILL_1_XOR2X1_14 INVX1_1/gnd DFFSR_53/S FILL
XFILL_0_NOR2X1_54 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_2_OAI21X1_2 BUFX2_79/A DFFSR_7/S FILL
XFILL_8_NAND3X1_142 INVX1_67/gnd DFFSR_175/S FILL
XINVX1_149 NOR3X1_5/A BUFX2_7/gnd INVX1_149/Y DFFSR_151/S INVX1
XFILL_1_1 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_12_DFFPOSX1_46 INVX1_39/gnd DFFSR_34/S FILL
XFILL_1_DFFSR_172 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_1_NAND2X1_123 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_15_XOR2X1_7 BUFX2_98/A DFFSR_6/S FILL
XFILL_42_DFFSR_203 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_7_AND2X2_13 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_46_DFFSR_94 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_18_DFFSR_102 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_5_DFFSR_279 BUFX2_99/A DFFSR_7/S FILL
XFILL_32_DFFSR_206 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_22_DFFSR_209 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_7_AND2X2_3 INVX1_1/gnd DFFSR_53/S FILL
XFILL_2_DFFSR_91 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_2_INVX1_38 AND2X2_38/B DFFSR_23/S FILL
XFILL_30_DFFSR_44 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_19_DFFSR_84 BUFX2_99/A DFFSR_7/S FILL
XFILL_12_DFFSR_212 OR2X2_2/gnd DFFSR_175/S FILL
XDFFSR_102 DFFSR_110/D DFFSR_45/CLK DFFSR_15/R DFFSR_98/S DFFSR_94/Q DFFSR_4/gnd DFFSR_98/S
+ DFFSR
XFILL_22_DFFPOSX1_35 INVX1_39/gnd DFFSR_54/S FILL
XFILL_15_CLKBUF1_7 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_6_NAND3X1_238 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_1_BUFX2_29 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_45_DFFSR_130 BUFX2_79/A DFFSR_6/S FILL
XFILL_8_DFFSR_206 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_35_DFFSR_133 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_49_DFFSR_237 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_25_DFFSR_136 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_39_DFFSR_240 INVX1_39/gnd DFFSR_34/S FILL
XFILL_1_INVX1_183 BUFX2_79/A DFFSR_6/S FILL
XFILL_27_DFFSR_91 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_38_DFFSR_51 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_49_DFFSR_11 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_1_CLKBUF1_4 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_7_NAND3X1_172 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_15_DFFSR_139 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_29_DFFSR_243 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_0_NAND2X1_153 BUFX2_98/A DFFSR_32/S FILL
XDFFSR_48 DFFSR_48/Q DFFSR_8/CLK DFFSR_8/R DFFSR_60/S DFFSR_40/Q DFFSR_8/gnd DFFSR_60/S
+ DFFSR
XFILL_19_DFFSR_246 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_11_DFFSR_41 BUFX2_98/A DFFSR_6/S FILL
XFILL_0_NOR2X1_18 OR2X2_4/gnd DFFSR_3/S FILL
XINVX1_113 DFFSR_216/Q BUFX2_77/gnd INVX1_113/Y DFFSR_98/S INVX1
XFILL_8_NAND3X1_106 INVX1_3/gnd DFFSR_23/S FILL
XFILL_12_DFFPOSX1_10 INVX1_67/gnd DFFSR_201/S FILL
XFILL_1_DFFSR_136 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_15_DFFSR_8 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_42_DFFSR_167 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_46_DFFSR_58 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_35_DFFSR_98 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_5_DFFSR_243 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_32_DFFSR_170 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_46_DFFSR_274 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_14_1_2 INVX1_39/gnd DFFSR_54/S FILL
XFILL_22_DFFSR_173 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_36_DFFSR_277 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_2_DFFSR_55 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_19_DFFSR_48 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_6_BUFX2_83 BUFX2_79/A DFFSR_7/S FILL
XFILL_12_DFFSR_176 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_4_AOI22X1_8 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_26_DFFSR_280 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_8_XOR2X1_12 INVX1_3/gnd DFFSR_23/S FILL
XFILL_20_CLKBUF1_38 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_6_NAND3X1_202 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_19_CLKBUF1_41 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_2_DFFPOSX1_21 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_36_DFFSR_4 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_8_DFFSR_170 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_49_DFFSR_201 INVX1_67/gnd DFFSR_201/S FILL
XAND2X2_17 NOR3X1_4/A NOR3X1_4/B XOR2X1_4/gnd BUFX2_34/A DFFSR_91/S AND2X2
XFILL_18_CLKBUF1_44 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_25_DFFSR_100 INVX1_1/gnd DFFSR_97/S FILL
XNAND3X1_238 INVX1_173/Y AOI21X1_36/B AOI21X1_36/A BUFX2_77/gnd NAND3X1_239/B DFFSR_98/S
+ NAND3X1
XFILL_39_DFFSR_204 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_17_CLKBUF1_47 BUFX2_98/A DFFSR_32/S FILL
XFILL_1_INVX1_147 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_38_DFFSR_15 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_27_DFFSR_55 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_16_DFFSR_95 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_4_AND2X2_14 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_15_DFFSR_103 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_2_DFFSR_280 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_7_NAND3X1_136 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_29_DFFSR_207 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_11_DFFPOSX1_40 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_0_NAND2X1_117 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_41_4_0 BUFX2_98/A DFFSR_32/S FILL
XDFFSR_12 DFFSR_68/D DFFSR_8/CLK DFFSR_8/R DFFSR_8/S DFFSR_12/D DFFSR_8/gnd DFFSR_8/S
+ DFFSR
XFILL_19_DFFSR_210 BUFX2_98/A DFFSR_6/S FILL
XFILL_39_6_1 BUFX2_79/A DFFSR_6/S FILL
XFILL_12_CLKBUF1_8 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_1_DFFSR_100 INVX1_1/gnd DFFSR_97/S FILL
XFILL_21_DFFPOSX1_29 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_42_DFFSR_131 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_46_DFFSR_22 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_35_DFFSR_62 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_5_DFFSR_207 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_32_DFFSR_134 INVX1_1/gnd DFFSR_53/S FILL
XFILL_46_DFFSR_238 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_5_NAND3X1_232 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_8_CLKBUF1_2 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_22_DFFSR_137 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_36_DFFSR_241 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_2_DFFSR_19 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_19_DFFSR_12 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_6_BUFX2_47 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_12_DFFSR_140 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_26_DFFSR_244 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_16_DFFSR_247 BUFX2_99/A DFFSR_7/S FILL
XFILL_45_2 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_6_NAND3X1_166 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_43_DFFSR_69 BUFX2_98/A DFFSR_32/S FILL
XFILL_8_DFFSR_134 INVX1_1/gnd DFFSR_53/S FILL
XFILL_49_DFFSR_165 BUFX2_72/gnd DFFSR_201/S FILL
XNAND3X1_202 INVX1_167/A INVX1_168/Y OAI21X1_78/C OR2X2_6/gnd NAND3X1_203/A DFFSR_53/S
+ NAND3X1
XFILL_39_DFFSR_168 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_17_CLKBUF1_11 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_27_DFFSR_19 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_16_DFFSR_59 AND2X2_38/B DFFSR_59/S FILL
XFILL_1_INVX1_111 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_7_NAND3X1_100 AND2X2_38/B DFFSR_59/S FILL
XFILL_2_DFFSR_244 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_3_BUFX2_94 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_29_DFFSR_171 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_16_CLKBUF1_14 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_43_DFFSR_275 BUFX2_99/A DFFSR_92/S FILL
XFILL_19_DFFSR_174 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_15_CLKBUF1_17 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_49_1_1 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_33_DFFSR_278 XOR2X1_1/gnd DFFSR_151/S FILL
XNOR2X1_56 NOR2X1_56/A NOR2X1_56/B AND2X2_38/B NOR2X1_56/Y DFFSR_59/S NOR2X1
XFILL_14_CLKBUF1_20 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_3_DFFSR_7 BUFX2_79/A DFFSR_7/S FILL
XFILL_1_AOI22X1_9 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_13_CLKBUF1_23 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_5_XOR2X1_13 INVX1_1/gnd DFFSR_97/S FILL
XFILL_4_NOR2X1_53 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_47_3_2 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_6_OAI21X1_1 BUFX2_79/A DFFSR_7/S FILL
XFILL_12_CLKBUF1_26 INVX1_1/gnd DFFSR_53/S FILL
XFILL_7_OAI21X1_118 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_7_DFFSR_73 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_24_DFFSR_66 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_35_DFFSR_26 BUFX2_79/A DFFSR_6/S FILL
XFILL_11_CLKBUF1_29 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_5_DFFSR_171 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_46_DFFSR_202 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_10_CLKBUF1_32 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_5_NAND3X1_196 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_22_DFFSR_101 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_9_DFFSR_278 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_36_DFFSR_205 INVX1_3/gnd DFFSR_79/S FILL
XFILL_1_DFFPOSX1_15 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_1_AND2X2_15 INVX1_3/gnd DFFSR_23/S FILL
XFILL_12_DFFSR_104 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_6_BUFX2_11 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_9_CLKBUF1_35 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_26_DFFSR_208 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_16_DFFSR_211 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_8_CLKBUF1_38 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_15_2_0 INVX1_39/gnd DFFSR_34/S FILL
XFILL_6_NAND3X1_130 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_7_CLKBUF1_41 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_10_DFFPOSX1_34 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_19_CLKBUF1_6 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_4_INVX1_67 INVX1_67/gnd DFFSR_201/S FILL
XFILL_43_DFFSR_33 BUFX2_98/A DFFSR_32/S FILL
XFILL_32_DFFSR_73 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_6_CLKBUF1_44 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_49_DFFSR_129 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_13_4_1 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_5_CLKBUF1_47 BUFX2_98/A DFFSR_32/S FILL
XNAND3X1_166 AOI22X1_20/D AOI22X1_20/C AOI21X1_15/Y DFFSR_34/gnd NAND3X1_167/B DFFSR_34/S
+ NAND3X1
XFILL_39_DFFSR_132 INVX1_3/gnd DFFSR_79/S FILL
XFILL_16_DFFSR_23 AND2X2_38/B DFFSR_23/S FILL
XCLKBUF1_44 clk DFFSR_1/gnd CLKBUF1_44/Y DFFSR_81/S CLKBUF1
XFILL_2_DFFSR_208 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_3_BUFX2_58 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_29_DFFSR_135 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_43_DFFSR_239 INVX1_39/gnd DFFSR_54/S FILL
XFILL_11_6_2 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_20_DFFPOSX1_23 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_5_CLKBUF1_3 BUFX2_98/A DFFSR_6/S FILL
XFILL_19_DFFSR_138 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_7_NOR3X1_4 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_33_DFFSR_242 OR2X2_3/gnd DFFSR_60/S FILL
XNOR2X1_20 NOR2X1_20/A NOR2X1_20/B OR2X2_4/gnd NOR2X1_20/Y DFFSR_32/S NOR2X1
XFILL_48_DFFSR_7 BUFX2_79/A DFFSR_7/S FILL
XFILL_4_NAND3X1_226 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_23_DFFSR_245 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_40_DFFSR_80 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_4_NOR2X1_17 BUFX2_79/A DFFSR_6/S FILL
XFILL_13_DFFSR_248 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_0_DFFPOSX1_45 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_7_DFFSR_37 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_50_7 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_13_DFFSR_70 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_24_DFFSR_30 BUFX2_98/A DFFSR_32/S FILL
XFILL_5_DFFSR_135 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_46_DFFSR_166 AND2X2_38/B DFFSR_59/S FILL
XFILL_5_NAND3X1_160 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_9_DFFSR_242 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_36_DFFSR_169 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_3_INVX1_9 BUFX2_99/A DFFSR_7/S FILL
XFILL_50_DFFSR_273 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_0_XOR2X1_7 BUFX2_98/A DFFSR_6/S FILL
XFILL_26_DFFSR_172 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_40_DFFSR_276 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_48_DFFSR_87 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_16_DFFSR_175 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_8_AOI22X1_7 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_30_DFFSR_279 BUFX2_99/A DFFSR_7/S FILL
XFILL_32_DFFSR_37 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_4_DFFSR_84 BUFX2_99/A DFFSR_7/S FILL
XFILL_4_INVX1_31 INVX1_1/gnd DFFSR_53/S FILL
XFILL_21_DFFSR_77 BUFX2_98/A DFFSR_32/S FILL
XFILL_2_XOR2X1_14 INVX1_1/gnd DFFSR_53/S FILL
XFILL_1_NOR2X1_54 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_3_OAI21X1_2 BUFX2_79/A DFFSR_7/S FILL
XFILL_5_CLKBUF1_11 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_21_1_2 BUFX2_8/gnd DFFSR_51/S FILL
XNAND3X1_130 INVX1_121/Y INVX1_122/Y INVX1_123/Y DFFSR_34/gnd NOR2X1_60/B DFFSR_34/S
+ NAND3X1
XFILL_4_CLKBUF1_14 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_2_DFFSR_172 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_3_BUFX2_22 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_3_0_1 INVX1_67/gnd DFFSR_175/S FILL
XFILL_43_DFFSR_203 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_3_CLKBUF1_17 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_8_AND2X2_13 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_19_DFFSR_102 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_6_DFFSR_279 BUFX2_99/A DFFSR_7/S FILL
XFILL_6_OAI21X1_112 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_33_DFFSR_206 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_14_DFFSR_5 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_13_NOR3X1_1 INVX1_3/gnd DFFSR_79/S FILL
XFILL_2_CLKBUF1_20 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_1_2_2 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_23_DFFSR_209 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_4_NAND3X1_190 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_1_CLKBUF1_23 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_40_DFFSR_44 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_29_DFFSR_84 BUFX2_99/A DFFSR_7/S FILL
XFILL_1_INVX1_78 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_13_DFFSR_212 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_0_CLKBUF1_26 INVX1_1/gnd DFFSR_53/S FILL
XFILL_16_CLKBUF1_7 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_13_DFFSR_34 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_0_BUFX2_69 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_46_DFFSR_130 BUFX2_79/A DFFSR_6/S FILL
XFILL_5_NAND3X1_124 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_9_DFFSR_206 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_36_DFFSR_133 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_48_4_0 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_50_DFFSR_237 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_26_DFFSR_136 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_35_DFFSR_1 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_10_4 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_40_DFFSR_240 INVX1_39/gnd DFFSR_34/S FILL
XFILL_2_INVX1_183 BUFX2_79/A DFFSR_6/S FILL
XFILL_37_DFFSR_91 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_48_DFFSR_51 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_2_CLKBUF1_4 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_16_DFFSR_139 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_46_6_1 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_30_DFFSR_243 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_20_DFFSR_246 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_4_DFFSR_48 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_21_DFFSR_41 BUFX2_98/A DFFSR_6/S FILL
XFILL_19_DFFPOSX1_17 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_10_DFFSR_81 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_1_NOR2X1_18 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_10_DFFSR_249 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_3_NAND3X1_220 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_2_DFFSR_136 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_27_DFFPOSX1_5 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_43_DFFSR_167 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_45_DFFSR_98 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_6_DFFSR_243 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_26_DFFPOSX1_8 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_33_DFFSR_170 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_47_DFFSR_274 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_4_NAND3X1_154 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_6_AND2X2_7 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_23_DFFSR_173 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_37_DFFSR_277 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_29_DFFSR_48 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_18_DFFSR_88 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_1_DFFSR_95 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_1_INVX1_42 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_13_DFFSR_176 OR2X2_6/gnd DFFSR_53/S FILL
XOAI21X1_112 NOR2X1_77/A XOR2X1_9/Y INVX1_212/Y BUFX2_8/gnd OR2X2_5/B DFFSR_81/S OAI21X1
XFILL_9_DFFPOSX1_28 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_5_AOI22X1_8 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_27_DFFSR_280 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_9_XOR2X1_12 INVX1_3/gnd DFFSR_23/S FILL
XFILL_0_BUFX2_33 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_0_OAI21X1_3 BUFX2_99/A DFFSR_92/S FILL
XFILL_9_DFFSR_170 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_50_DFFSR_201 INVX1_67/gnd DFFSR_201/S FILL
XFILL_18_DFFPOSX1_47 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_26_DFFSR_100 INVX1_1/gnd DFFSR_97/S FILL
XFILL_40_DFFSR_204 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_2_INVX1_147 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_48_DFFSR_15 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_37_DFFSR_55 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_26_DFFSR_95 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_5_AND2X2_14 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_16_DFFSR_103 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_3_DFFSR_280 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_30_DFFSR_207 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_54_3_2 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_20_DFFSR_210 BUFX2_98/A DFFSR_6/S FILL
XFILL_4_DFFSR_12 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_10_DFFSR_45 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_5_OAI21X1_106 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_10_DFFSR_213 INVX1_3/gnd DFFSR_23/S FILL
XFILL_3_NAND3X1_184 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_13_CLKBUF1_8 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_2_DFFSR_4 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_2_DFFSR_100 INVX1_1/gnd DFFSR_97/S FILL
XFILL_43_DFFSR_131 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_45_DFFSR_62 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_6_DFFSR_207 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_33_DFFSR_134 INVX1_1/gnd DFFSR_53/S FILL
XFILL_47_DFFSR_238 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_22_2_0 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_9_CLKBUF1_2 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_23_DFFSR_137 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_4_NAND3X1_118 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_37_DFFSR_241 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_29_DFFSR_12 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_18_DFFSR_52 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_1_DFFSR_59 AND2X2_38/B DFFSR_59/S FILL
XFILL_5_BUFX2_87 INVX1_1/gnd DFFSR_53/S FILL
XFILL_13_DFFSR_140 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_27_DFFSR_244 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_6_NAND2X1_154 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_0_OR2X2_4 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_20_4_1 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_17_DFFSR_247 BUFX2_99/A DFFSR_7/S FILL
XFILL_2_3_0 INVX1_67/gnd DFFSR_201/S FILL
XFILL_26_DFFSR_8 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_9_DFFSR_134 INVX1_1/gnd DFFSR_53/S FILL
XFILL_18_6_2 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_18_DFFPOSX1_11 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_50_DFFSR_165 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_0_5_1 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_40_DFFSR_168 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_37_DFFSR_19 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_9_DFFSR_66 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_2_INVX1_111 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_15_DFFSR_99 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_26_DFFSR_59 AND2X2_38/B DFFSR_59/S FILL
XFILL_3_DFFSR_244 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_2_NAND3X1_214 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_30_DFFSR_171 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_44_DFFSR_275 BUFX2_99/A DFFSR_92/S FILL
XFILL_20_DFFSR_174 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_34_DFFSR_278 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_16_DFFPOSX1_2 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_10_DFFSR_177 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_2_AOI22X1_9 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_15_DFFPOSX1_5 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_6_XOR2X1_13 INVX1_1/gnd DFFSR_97/S FILL
XFILL_3_NAND3X1_148 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_5_NOR2X1_53 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_47_DFFSR_4 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_14_DFFPOSX1_8 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_7_OAI21X1_1 BUFX2_79/A DFFSR_7/S FILL
XFILL_8_DFFPOSX1_22 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_34_DFFSR_66 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_45_DFFSR_26 BUFX2_79/A DFFSR_6/S FILL
XFILL_6_DFFSR_171 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_47_DFFSR_202 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_23_DFFSR_101 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_37_DFFSR_205 INVX1_3/gnd DFFSR_79/S FILL
XFILL_18_DFFSR_16 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_1_DFFSR_23 AND2X2_38/B DFFSR_23/S FILL
XFILL_2_AND2X2_15 INVX1_3/gnd DFFSR_23/S FILL
XBUFX2_91 BUFX2_91/A DFFSR_28/gnd BUFX2_91/Y DFFSR_3/S BUFX2
XFILL_13_DFFSR_104 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_5_BUFX2_51 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_17_DFFPOSX1_41 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_27_DFFSR_208 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_6_NAND2X1_118 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_2_INVX1_6 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_17_DFFSR_211 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_28_1_2 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_1_NAND3X1_244 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_0_NOR2X1_4 INVX1_1/gnd DFFSR_53/S FILL
XFILL_20_CLKBUF1_6 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_42_DFFSR_73 OR2X2_1/gnd DFFSR_51/S FILL
XNAND2X1_154 NAND2X1_153/B INVX1_208/Y OR2X2_4/gnd AOI21X1_53/A DFFSR_3/S NAND2X1
XFILL_10_CLKBUF1_9 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_50_DFFSR_129 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_4_OAI21X1_100 INVX1_3/gnd DFFSR_79/S FILL
XFILL_8_AOI21X1_46 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_27_DFFPOSX1_30 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_40_DFFSR_132 INVX1_3/gnd DFFSR_79/S FILL
XFILL_7_AOI21X1_49 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_8_2_2 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_9_DFFSR_30 BUFX2_98/A DFFSR_32/S FILL
XFILL_15_DFFSR_63 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_2_NAND3X1_178 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_26_DFFSR_23 AND2X2_38/B DFFSR_23/S FILL
XFILL_3_DFFSR_208 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_2_BUFX2_98 BUFX2_79/A DFFSR_7/S FILL
XFILL_30_DFFSR_135 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_6_AOI21X1_52 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_44_DFFSR_239 INVX1_39/gnd DFFSR_54/S FILL
XFILL_6_CLKBUF1_3 BUFX2_98/A DFFSR_6/S FILL
XFILL_20_DFFSR_138 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_5_AOI21X1_55 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_34_DFFSR_242 OR2X2_3/gnd DFFSR_60/S FILL
XAOI21X1_52 AOI21X1_52/A AOI21X1_52/B NOR3X1_6/A OR2X2_6/gnd AOI21X1_52/Y DFFSR_53/S
+ AOI21X1
XFILL_10_DFFSR_141 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_4_AOI21X1_58 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_24_DFFSR_245 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_50_DFFSR_80 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_5_NOR2X1_17 BUFX2_79/A DFFSR_6/S FILL
XFILL_13_DFFSR_2 BUFX2_79/A DFFSR_7/S FILL
XFILL_3_NAND3X1_112 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_14_DFFSR_248 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_3_AOI21X1_61 AND2X2_38/B DFFSR_59/S FILL
XFILL_2_AOI21X1_64 AND2X2_38/B DFFSR_59/S FILL
XFILL_54_4 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_5_NAND2X1_148 INVX1_67/gnd DFFSR_175/S FILL
XFILL_23_DFFSR_70 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_34_DFFSR_30 BUFX2_98/A DFFSR_32/S FILL
XFILL_6_DFFSR_77 BUFX2_98/A DFFSR_32/S FILL
XFILL_1_AOI21X1_67 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_6_DFFSR_135 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_47_DFFSR_166 AND2X2_38/B DFFSR_59/S FILL
XFILL_0_AOI21X1_70 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_53_6_1 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_37_DFFSR_169 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_5_BUFX2_15 DFFSR_8/gnd DFFSR_8/S FILL
XBUFX2_55 BUFX2_53/A DFFSR_1/gnd BUFX2_55/Y DFFSR_1/S BUFX2
XFILL_0_DFFSR_245 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_27_DFFSR_172 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_41_DFFSR_276 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_17_DFFSR_175 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_8_OAI21X1_94 INVX1_67/gnd DFFSR_175/S FILL
XFILL_9_AOI22X1_7 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_31_DFFSR_279 BUFX2_99/A DFFSR_7/S FILL
XFILL_1_NAND3X1_208 DFFSR_46/gnd DFFSR_54/S FILL
XOAI21X1_5 INVX1_37/Y OAI21X1_4/B OAI21X1_5/C DFFSR_8/gnd NOR2X1_19/B DFFSR_8/S OAI21X1
XFILL_7_OAI21X1_97 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_42_DFFSR_37 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_3_INVX1_71 BUFX2_79/A DFFSR_6/S FILL
XFILL_31_DFFSR_77 BUFX2_98/A DFFSR_32/S FILL
XFILL_3_XOR2X1_14 INVX1_1/gnd DFFSR_53/S FILL
XNAND2X1_118 DFFSR_79/S din[2] NOR3X1_6/gnd OAI21X1_87/C DFFSR_79/S NAND2X1
XFILL_2_NOR2X1_54 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_4_OAI21X1_2 BUFX2_79/A DFFSR_7/S FILL
XFILL_8_AOI21X1_10 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_7_AOI21X1_13 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_2_NAND3X1_142 INVX1_67/gnd DFFSR_175/S FILL
XFILL_15_DFFSR_27 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_3_DFFSR_172 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_2_BUFX2_62 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_6_AOI21X1_16 INVX1_67/gnd DFFSR_175/S FILL
XFILL_44_DFFSR_203 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_9_AND2X2_13 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_7_DFFPOSX1_16 INVX1_67/gnd DFFSR_175/S FILL
XFILL_20_DFFSR_102 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_7_DFFSR_279 BUFX2_99/A DFFSR_7/S FILL
XFILL_4_NAND2X1_178 INVX1_1/gnd DFFSR_53/S FILL
XFILL_4_DFFPOSX1_2 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_5_AOI21X1_19 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_34_DFFSR_206 OR2X2_2/gnd DFFSR_175/S FILL
XAOI21X1_16 INVX1_153/Y INVX1_140/A INVX1_141/Y INVX1_67/gnd AOI21X1_16/Y DFFSR_175/S
+ AOI21X1
XFILL_10_DFFSR_105 INVX1_1/gnd DFFSR_53/S FILL
XFILL_3_DFFPOSX1_5 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_4_AOI21X1_22 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_24_DFFSR_209 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_50_DFFSR_44 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_39_DFFSR_84 BUFX2_99/A DFFSR_7/S FILL
XFILL_2_DFFPOSX1_8 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_3_AOI21X1_25 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_14_DFFSR_212 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_2_AOI21X1_28 AND2X2_38/B DFFSR_23/S FILL
XFILL_16_DFFPOSX1_35 INVX1_39/gnd DFFSR_54/S FILL
XFILL_5_NAND2X1_112 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_17_CLKBUF1_7 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_6_DFFSR_41 BUFX2_98/A DFFSR_6/S FILL
XFILL_23_DFFSR_34 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_12_DFFSR_74 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_1_AOI21X1_31 INVX1_39/gnd DFFSR_34/S FILL
XFILL_0_NAND3X1_238 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_47_DFFSR_130 BUFX2_79/A DFFSR_6/S FILL
XFILL_0_AOI21X1_34 INVX1_39/gnd DFFSR_34/S FILL
XFILL_37_DFFSR_133 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_0_DFFSR_209 BUFX2_72/gnd DFFSR_276/S FILL
XBUFX2_19 AND2X2_4/Y DFFSR_28/gnd BUFX2_19/Y DFFSR_3/S BUFX2
XFILL_14_1 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_27_DFFSR_136 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_26_DFFPOSX1_24 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_3_INVX1_183 BUFX2_79/A DFFSR_6/S FILL
XFILL_41_DFFSR_240 INVX1_39/gnd DFFSR_34/S FILL
XFILL_47_DFFSR_91 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_3_CLKBUF1_4 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_17_DFFSR_139 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_8_OAI21X1_58 INVX1_39/gnd DFFSR_54/S FILL
XFILL_31_DFFSR_243 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_1_NAND3X1_172 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_6_NAND2X1_79 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_7_OAI21X1_61 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_21_DFFSR_246 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_3_INVX1_35 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_3_DFFSR_88 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_31_DFFSR_41 BUFX2_98/A DFFSR_6/S FILL
XFILL_20_DFFSR_81 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_2_NOR2X1_18 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_6_DFFPOSX1_46 INVX1_39/gnd DFFSR_34/S FILL
XFILL_11_DFFSR_249 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_6_OAI21X1_64 INVX1_1/gnd DFFSR_53/S FILL
XFILL_5_NAND2X1_82 DFFSR_1/gnd DFFSR_81/S FILL
XNAND2X1_79 OAI21X1_42/Y NAND2X1_79/B XOR2X1_1/gnd NAND2X1_79/Y DFFSR_151/S NAND2X1
XFILL_5_OAI21X1_67 INVX1_1/gnd DFFSR_97/S FILL
XFILL_4_NAND2X1_85 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_29_2_0 NOR3X1_6/gnd DFFSR_91/S FILL
XOAI21X1_64 INVX1_134/Y NOR2X1_69/B OAI21X1_63/Y INVX1_1/gnd AOI22X1_26/B DFFSR_53/S
+ OAI21X1
XFILL_2_NAND3X1_106 INVX1_3/gnd DFFSR_23/S FILL
XFILL_3_DFFSR_136 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_4_OAI21X1_70 INVX1_3/gnd DFFSR_23/S FILL
XFILL_3_NAND2X1_88 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_2_BUFX2_26 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_44_DFFSR_167 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_2_NAND2X1_91 INVX1_39/gnd DFFSR_54/S FILL
XFILL_3_OAI21X1_73 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_7_DFFSR_243 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_1_DFFSR_1 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_4_NAND2X1_142 INVX1_67/gnd DFFSR_175/S FILL
XFILL_34_DFFSR_170 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_27_4_1 INVX1_3/gnd DFFSR_79/S FILL
XFILL_48_DFFSR_274 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_12_NOR3X1_5 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_1_NAND2X1_94 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_2_OAI21X1_76 INVX1_1/gnd DFFSR_53/S FILL
XFILL_24_DFFSR_173 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_1_OAI21X1_79 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_0_NAND2X1_97 INVX1_1/gnd DFFSR_97/S FILL
XFILL_9_3_0 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_38_DFFSR_277 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_0_INVX1_82 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_39_DFFSR_48 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_28_DFFSR_88 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_14_DFFSR_176 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_0_OAI21X1_82 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_25_6_2 AND2X2_38/B DFFSR_23/S FILL
XFILL_6_AOI22X1_8 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_28_DFFSR_280 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_7_5_1 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_12_DFFSR_38 BUFX2_98/A DFFSR_6/S FILL
XFILL_0_XOR2X1_15 BUFX2_99/A DFFSR_7/S FILL
XFILL_1_OAI21X1_3 BUFX2_99/A DFFSR_92/S FILL
XFILL_0_NAND3X1_202 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_0_DFFSR_173 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_25_DFFSR_5 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_27_DFFSR_100 INVX1_1/gnd DFFSR_97/S FILL
XFILL_41_DFFSR_204 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_3_INVX1_147 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_47_DFFSR_55 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_36_DFFSR_95 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_6_AND2X2_14 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_17_DFFSR_103 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_4_DFFSR_280 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_8_OAI21X1_22 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_1_NAND3X1_136 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_31_DFFSR_207 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_6_NAND2X1_43 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_21_DFFSR_210 BUFX2_98/A DFFSR_6/S FILL
XFILL_7_OAI21X1_25 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_3_DFFSR_52 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_20_DFFSR_45 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_6_DFFPOSX1_10 INVX1_67/gnd DFFSR_201/S FILL
XFILL_6_OAI21X1_28 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_11_DFFSR_213 INVX1_3/gnd DFFSR_23/S FILL
XFILL_3_NAND2X1_172 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_5_NAND2X1_46 INVX1_39/gnd DFFSR_34/S FILL
XNAND2X1_43 DFFSR_236/Q NOR2X1_34/Y BUFX2_8/gnd NAND2X1_43/Y DFFSR_81/S NAND2X1
XFILL_4_NAND2X1_49 INVX1_3/gnd DFFSR_79/S FILL
XFILL_5_OAI21X1_31 AND2X2_38/B DFFSR_23/S FILL
XFILL_14_CLKBUF1_8 NOR3X1_6/gnd DFFSR_79/S FILL
XOAI21X1_28 INVX1_131/Y NAND2X1_65/Y OAI21X1_27/Y XOR2X1_1/gnd OAI21X1_28/Y DFFSR_151/S
+ OAI21X1
XFILL_4_OAI21X1_34 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_3_NAND2X1_52 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_3_DFFSR_100 INVX1_1/gnd DFFSR_97/S FILL
XDFFPOSX1_46 AND2X2_34/B CLKBUF1_49/Y NOR2X1_79/Y INVX1_39/gnd DFFSR_34/S DFFPOSX1
XFILL_44_DFFSR_131 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_2_NAND2X1_55 INVX1_39/gnd DFFSR_34/S FILL
XFILL_15_DFFPOSX1_29 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_3_OAI21X1_37 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_46_DFFSR_1 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_7_DFFSR_207 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_4_NAND2X1_106 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_34_DFFSR_134 INVX1_1/gnd DFFSR_53/S FILL
XFILL_48_DFFSR_238 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_1_NAND2X1_58 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_2_OAI21X1_40 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_35_1_2 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_24_DFFSR_137 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_0_NAND2X1_61 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_1_OAI21X1_43 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_38_DFFSR_241 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_39_DFFSR_12 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_28_DFFSR_52 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_0_INVX1_46 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_0_INVX1_184 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_0_DFFSR_99 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_17_DFFSR_92 BUFX2_99/A DFFSR_92/S FILL
XFILL_0_CLKBUF1_5 BUFX2_99/A DFFSR_92/S FILL
XFILL_19_6 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_14_DFFSR_140 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_0_OAI21X1_46 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_28_DFFSR_244 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_36_1 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_18_DFFSR_247 BUFX2_99/A DFFSR_7/S FILL
XFILL_25_DFFPOSX1_18 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_9_AOI22X1_12 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_1_INVX1_3 INVX1_3/gnd DFFSR_79/S FILL
XFILL_0_NAND3X1_166 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_8_AOI22X1_15 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_7_AOI22X1_18 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_5_DFFPOSX1_40 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_0_DFFSR_137 BUFX2_7/gnd DFFSR_216/S FILL
XDFFSR_247 INVX1_110/A CLKBUF1_3/Y BUFX2_65/Y DFFSR_7/S DFFSR_239/Q BUFX2_99/A DFFSR_7/S
+ DFFSR
XFILL_6_AOI22X1_21 AND2X2_38/B DFFSR_59/S FILL
XFILL_41_DFFSR_168 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_47_DFFSR_19 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_3_INVX1_111 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_25_DFFSR_99 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_36_DFFSR_59 AND2X2_38/B DFFSR_59/S FILL
XFILL_4_DFFSR_244 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_5_AOI22X1_24 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_1_NAND3X1_100 AND2X2_38/B DFFSR_59/S FILL
XFILL_31_DFFSR_171 BUFX2_8/gnd DFFSR_81/S FILL
XAOI22X1_21 AND2X2_32/Y AND2X2_33/Y AOI22X1_21/C INVX1_151/Y AND2X2_38/B AOI21X1_27/C
+ DFFSR_59/S AOI22X1
XFILL_45_DFFSR_275 BUFX2_99/A DFFSR_92/S FILL
XFILL_4_AOI22X1_27 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_21_DFFSR_174 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_3_DFFSR_16 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_35_DFFSR_278 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_3_NAND2X1_136 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_5_NAND2X1_10 BUFX2_79/A DFFSR_7/S FILL
XFILL_11_DFFSR_177 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_3_AOI22X1_9 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_4_NAND2X1_13 BUFX2_99/A DFFSR_92/S FILL
XFILL_7_XOR2X1_13 INVX1_1/gnd DFFSR_97/S FILL
XFILL_6_NOR2X1_53 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_8_OAI21X1_1 BUFX2_79/A DFFSR_7/S FILL
XFILL_3_NAND2X1_16 BUFX2_79/A DFFSR_7/S FILL
XDFFPOSX1_10 BUFX2_7/A CLKBUF1_43/Y NOR2X1_62/Y INVX1_67/gnd DFFSR_201/S DFFPOSX1
XFILL_2_NAND2X1_19 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_44_DFFSR_66 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_1_OAI21X1_118 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_7_DFFSR_171 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_24_DFFPOSX1_48 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_1_NAND2X1_22 BUFX2_99/A DFFSR_7/S FILL
XFILL_48_DFFSR_202 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_24_DFFSR_101 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_8_NAND3X1_78 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_0_NAND2X1_25 BUFX2_99/A DFFSR_7/S FILL
XFILL_0_INVX1_148 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_28_DFFSR_16 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_0_DFFSR_63 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_0_INVX1_10 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_38_DFFSR_205 INVX1_3/gnd DFFSR_79/S FILL
XFILL_17_DFFSR_56 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_3_AND2X2_15 INVX1_3/gnd DFFSR_23/S FILL
XFILL_14_DFFSR_104 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_7_NAND3X1_81 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_4_BUFX2_91 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_0_OAI21X1_10 BUFX2_79/A DFFSR_7/S FILL
XFILL_28_DFFSR_208 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_6_NAND3X1_84 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_18_DFFSR_211 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_5_NAND3X1_87 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_0_NAND3X1_130 DFFSR_34/gnd DFFSR_34/S FILL
XNAND3X1_84 NAND3X1_84/A NAND3X1_84/B AND2X2_21/Y DFFSR_34/gnd NOR2X1_43/A DFFSR_34/S
+ NAND3X1
XFILL_4_NAND3X1_90 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_11_CLKBUF1_9 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_3_NAND3X1_93 XOR2X1_1/gnd DFFSR_208/S FILL
XDFFSR_211 INVX1_78/A CLKBUF1_11/Y BUFX2_68/Y DFFSR_216/S INVX1_79/A BUFX2_7/gnd DFFSR_216/S
+ DFFSR
XFILL_0_DFFSR_101 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_2_NAND2X1_166 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_41_DFFSR_132 INVX1_3/gnd DFFSR_79/S FILL
XFILL_2_NAND3X1_96 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_8_DFFSR_70 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_25_DFFSR_63 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_36_DFFSR_23 AND2X2_38/B DFFSR_23/S FILL
XFILL_4_DFFSR_208 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_1_NAND3X1_99 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_31_DFFSR_135 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_45_DFFSR_239 INVX1_39/gnd DFFSR_54/S FILL
XFILL_7_CLKBUF1_3 BUFX2_98/A DFFSR_6/S FILL
XFILL_21_DFFSR_138 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_14_DFFPOSX1_23 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_35_DFFSR_242 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_11_DFFSR_141 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_3_NAND2X1_100 INVX1_39/gnd DFFSR_54/S FILL
XFILL_25_DFFSR_245 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_6_NOR2X1_17 BUFX2_79/A DFFSR_6/S FILL
XFILL_15_DFFSR_248 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_11_OAI22X1_18 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_37_DFFSR_8 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_10_OAI22X1_21 BUFX2_98/A DFFSR_32/S FILL
XFILL_44_DFFSR_30 BUFX2_98/A DFFSR_32/S FILL
XFILL_33_DFFSR_70 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_7_DFFSR_135 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_24_DFFPOSX1_12 AND2X2_38/B DFFSR_23/S FILL
XFILL_9_NAND3X1_39 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_48_DFFSR_166 AND2X2_38/B DFFSR_59/S FILL
XFILL_9_OAI22X1_24 BUFX2_98/A DFFSR_32/S FILL
XFILL_8_NAND3X1_42 BUFX2_79/A DFFSR_6/S FILL
XFILL_0_DFFSR_27 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_0_INVX1_112 AND2X2_38/B DFFSR_23/S FILL
XFILL_8_NAND3X1_215 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_38_DFFSR_169 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_17_DFFSR_20 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_8_OAI22X1_27 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_7_NAND3X1_45 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_1_DFFSR_245 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_4_BUFX2_55 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_4_DFFPOSX1_34 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_28_DFFSR_172 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_42_DFFSR_276 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_6_NAND3X1_48 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_7_OAI22X1_30 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_18_DFFSR_175 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_32_DFFSR_279 BUFX2_99/A DFFSR_7/S FILL
XFILL_8_NOR3X1_1 INVX1_3/gnd DFFSR_79/S FILL
XFILL_5_NAND3X1_51 BUFX2_99/A DFFSR_7/S FILL
XFILL_6_OAI22X1_33 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_36_2_0 BUFX2_99/A DFFSR_92/S FILL
XNAND3X1_48 NOR2X1_21/Y NOR2X1_22/Y NOR2X1_23/Y OR2X2_4/gnd XOR2X1_14/A DFFSR_3/S
+ NAND3X1
XFILL_5_OAI22X1_36 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_4_NAND3X1_54 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_41_DFFSR_77 BUFX2_98/A DFFSR_32/S FILL
XFILL_4_XOR2X1_14 INVX1_1/gnd DFFSR_53/S FILL
XFILL_3_NOR2X1_54 BUFX2_8/gnd DFFSR_51/S FILL
XOAI22X1_33 INVX1_80/Y OAI22X1_45/B INVX1_81/Y OAI22X1_45/D OR2X2_1/gnd NOR2X1_42/A
+ DFFSR_51/S OAI22X1
XFILL_3_NAND3X1_57 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_5_OAI21X1_2 BUFX2_79/A DFFSR_7/S FILL
XDFFSR_175 DFFSR_191/D CLKBUF1_10/Y BUFX2_64/Y DFFSR_175/S DFFSR_175/D OR2X2_2/gnd
+ DFFSR_175/S DFFSR
XFILL_4_OAI22X1_39 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_34_4_1 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_2_NAND2X1_130 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_2_NAND3X1_60 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_3_OAI22X1_42 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_8_DFFSR_34 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_25_DFFSR_27 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_14_DFFSR_67 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_4_DFFSR_172 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_2_OAI22X1_45 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_1_NAND3X1_63 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_32_6_2 INVX1_1/gnd DFFSR_97/S FILL
XFILL_45_DFFSR_203 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_0_NAND3X1_66 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_21_DFFSR_102 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_8_DFFSR_279 BUFX2_99/A DFFSR_7/S FILL
XFILL_1_OAI22X1_48 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_35_DFFSR_206 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_0_OAI21X1_112 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_0_AND2X2_16 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_11_DFFSR_105 INVX1_1/gnd DFFSR_53/S FILL
XFILL_23_DFFPOSX1_42 INVX1_39/gnd DFFSR_34/S FILL
XFILL_0_OAI22X1_51 INVX1_39/gnd DFFSR_54/S FILL
XFILL_25_DFFSR_209 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_1_XOR2X1_4 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_49_DFFSR_84 BUFX2_99/A DFFSR_7/S FILL
XFILL_15_DFFSR_212 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_7_NAND3X1_245 OR2X2_4/gnd DFFSR_3/S FILL
XINVX1_68 INVX1_68/A INVX1_67/gnd INVX1_68/Y DFFSR_201/S INVX1
XFILL_18_CLKBUF1_7 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_5_DFFSR_81 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_33_DFFSR_34 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_22_DFFSR_74 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_48_DFFSR_130 BUFX2_79/A DFFSR_6/S FILL
XFILL_38_DFFSR_133 BUFX2_77/gnd DFFSR_5/S FILL
XINVX1_186 DFFSR_6/D BUFX2_79/A INVX1_186/Y DFFSR_6/S INVX1
XFILL_8_NAND3X1_179 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_1_DFFSR_209 BUFX2_72/gnd DFFSR_276/S FILL
XCLKBUF1_7 BUFX2_6/Y OR2X2_4/gnd CLKBUF1_7/Y DFFSR_32/S CLKBUF1
XFILL_4_BUFX2_19 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_28_DFFSR_136 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_1_NAND2X1_160 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_4_INVX1_183 BUFX2_79/A DFFSR_6/S FILL
XFILL_42_DFFSR_240 INVX1_39/gnd DFFSR_34/S FILL
XFILL_6_NAND3X1_12 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_4_CLKBUF1_4 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_18_DFFSR_139 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_32_DFFSR_243 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_24_DFFSR_2 BUFX2_79/A DFFSR_7/S FILL
XFILL_5_NAND3X1_15 DFFSR_4/gnd DFFSR_4/S FILL
XNAND3X1_12 NAND2X1_14/Y NAND3X1_9/Y AND2X2_7/Y OR2X2_4/gnd NOR2X1_11/A DFFSR_32/S
+ NAND3X1
XFILL_22_DFFSR_246 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_4_NAND3X1_18 BUFX2_79/A DFFSR_7/S FILL
XFILL_41_DFFSR_41 BUFX2_98/A DFFSR_6/S FILL
XFILL_2_INVX1_75 BUFX2_98/A DFFSR_6/S FILL
XFILL_30_DFFSR_81 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_3_NOR2X1_18 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_13_DFFPOSX1_17 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_12_DFFSR_249 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_3_NAND3X1_21 OR2X2_6/gnd DFFSR_53/S FILL
XDFFSR_139 DFFSR_195/D CLKBUF1_17/Y BUFX2_69/Y DFFSR_34/S INVX1_76/A DFFSR_34/gnd
+ DFFSR_34/S DFFSR
XFILL_42_1_2 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_2_NAND3X1_24 INVX1_1/gnd DFFSR_97/S FILL
XFILL_14_DFFSR_31 BUFX2_79/A DFFSR_6/S FILL
XFILL_4_DFFSR_136 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_1_NAND3X1_27 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_1_BUFX2_66 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_45_DFFSR_167 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_8_DFFSR_243 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_1_OAI22X1_12 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_0_NAND3X1_30 BUFX2_79/A DFFSR_6/S FILL
XFILL_35_DFFSR_170 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_49_DFFSR_274 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_0_OAI22X1_15 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_25_DFFSR_173 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_39_DFFSR_277 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_49_DFFSR_48 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_38_DFFSR_88 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_15_DFFSR_176 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_7_NAND3X1_209 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_7_AOI22X1_8 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_29_DFFSR_280 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_3_DFFPOSX1_28 BUFX2_72/gnd DFFSR_201/S FILL
XDFFSR_85 INVX1_33/A DFFSR_85/CLK DFFSR_3/R DFFSR_8/S DFFSR_77/Q DFFSR_8/gnd DFFSR_8/S
+ DFFSR
XINVX1_32 INVX1_32/A OR2X2_6/gnd INVX1_32/Y DFFSR_53/S INVX1
XFILL_5_DFFSR_45 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_10_0_0 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_11_DFFSR_78 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_22_DFFSR_38 BUFX2_98/A DFFSR_6/S FILL
XFILL_1_XOR2X1_15 BUFX2_99/A DFFSR_7/S FILL
XFILL_0_NOR2X1_55 INVX1_39/gnd DFFSR_54/S FILL
XFILL_2_OAI21X1_3 BUFX2_99/A DFFSR_92/S FILL
XFILL_8_NAND3X1_143 BUFX2_8/gnd DFFSR_51/S FILL
XINVX1_150 AND2X2_35/B BUFX2_8/gnd INVX1_150/Y DFFSR_81/S INVX1
XFILL_1_DFFSR_173 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_1_2 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_12_DFFPOSX1_47 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_28_DFFSR_100 INVX1_1/gnd DFFSR_97/S FILL
XFILL_1_NAND2X1_124 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_15_XOR2X1_8 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_42_DFFSR_204 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_4_INVX1_147 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_46_DFFSR_95 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_7_AND2X2_14 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_18_DFFSR_103 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_5_DFFSR_280 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_32_DFFSR_207 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_22_DFFSR_210 BUFX2_98/A DFFSR_6/S FILL
XFILL_7_AND2X2_4 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_19_DFFSR_85 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_30_DFFSR_45 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_2_DFFSR_92 BUFX2_99/A DFFSR_92/S FILL
XFILL_2_INVX1_39 INVX1_39/gnd DFFSR_34/S FILL
XFILL_12_DFFSR_213 INVX1_3/gnd DFFSR_23/S FILL
XFILL_22_DFFPOSX1_36 OR2X2_2/gnd DFFSR_175/S FILL
XDFFSR_103 AOI22X1_7/B CLKBUF1_5/Y DFFSR_9/R DFFSR_60/S DFFSR_95/Q DFFSR_8/gnd DFFSR_60/S
+ DFFSR
XFILL_15_CLKBUF1_8 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_4_DFFSR_100 INVX1_1/gnd DFFSR_97/S FILL
XFILL_6_NAND3X1_239 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_1_BUFX2_30 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_45_DFFSR_131 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_8_DFFSR_207 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_35_DFFSR_134 INVX1_1/gnd DFFSR_53/S FILL
XFILL_49_DFFSR_238 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_25_DFFSR_137 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_39_DFFSR_241 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_49_DFFSR_12 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_1_INVX1_184 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_38_DFFSR_52 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_27_DFFSR_92 BUFX2_99/A DFFSR_92/S FILL
XFILL_1_CLKBUF1_5 BUFX2_99/A DFFSR_92/S FILL
XFILL_15_DFFSR_140 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_7_NAND3X1_173 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_29_DFFSR_244 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_0_NAND2X1_154 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_19_DFFSR_247 BUFX2_99/A DFFSR_7/S FILL
XDFFSR_49 INVX1_1/A DFFSR_9/CLK BUFX2_49/Y DFFSR_92/S INVX1_2/A OR2X2_6/gnd DFFSR_92/S
+ DFFSR
XFILL_11_DFFSR_42 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_0_NOR2X1_19 DFFSR_28/gnd DFFSR_3/S FILL
XINVX1_114 DFFSR_216/D BUFX2_77/gnd INVX1_114/Y DFFSR_98/S INVX1
XFILL_8_NAND3X1_107 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_1_DFFSR_137 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_12_DFFPOSX1_11 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_15_DFFSR_9 BUFX2_79/A DFFSR_6/S FILL
XFILL_42_DFFSR_168 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_4_INVX1_111 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_35_DFFSR_99 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_46_DFFSR_59 AND2X2_38/B DFFSR_59/S FILL
XFILL_5_DFFSR_244 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_32_DFFSR_171 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_46_DFFSR_275 BUFX2_99/A DFFSR_92/S FILL
XFILL_22_DFFSR_174 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_2_DFFSR_56 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_19_DFFSR_49 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_36_DFFSR_278 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_12_DFFSR_177 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_6_BUFX2_84 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_4_AOI22X1_9 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_8_XOR2X1_13 INVX1_1/gnd DFFSR_97/S FILL
XFILL_9_OAI21X1_1 BUFX2_79/A DFFSR_7/S FILL
XFILL_20_CLKBUF1_39 INVX1_1/gnd DFFSR_53/S FILL
XFILL_6_NAND3X1_203 INVX1_1/gnd DFFSR_97/S FILL
XFILL_19_CLKBUF1_42 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_36_DFFSR_5 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_2_DFFPOSX1_22 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_8_DFFSR_171 BUFX2_8/gnd DFFSR_81/S FILL
XAND2X2_18 BUFX2_32/Y AND2X2_18/B AND2X2_38/B AND2X2_18/Y DFFSR_59/S AND2X2
XFILL_18_CLKBUF1_45 BUFX2_79/A DFFSR_7/S FILL
XFILL_49_DFFSR_202 NOR3X1_6/gnd DFFSR_91/S FILL
XNAND3X1_239 NAND3X1_239/A NAND3X1_239/B INVX1_179/Y DFFSR_8/gnd AOI21X1_38/A DFFSR_60/S
+ NAND3X1
XFILL_25_DFFSR_101 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_43_2_0 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_1_INVX1_148 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_38_DFFSR_16 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_17_CLKBUF1_48 INVX1_3/gnd DFFSR_79/S FILL
XFILL_39_DFFSR_205 INVX1_3/gnd DFFSR_79/S FILL
XFILL_27_DFFSR_56 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_16_DFFSR_96 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_4_AND2X2_15 INVX1_3/gnd DFFSR_23/S FILL
XFILL_7_NAND3X1_137 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_15_DFFSR_104 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_29_DFFSR_208 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_11_DFFPOSX1_41 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_19_DFFSR_211 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_41_4_1 BUFX2_98/A DFFSR_32/S FILL
XDFFSR_13 DFFSR_13/Q DFFSR_9/CLK DFFSR_73/R DFFSR_53/S INVX1_31/A OR2X2_6/gnd DFFSR_53/S
+ DFFSR
XFILL_0_NAND2X1_118 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_39_6_2 BUFX2_79/A DFFSR_6/S FILL
XFILL_12_CLKBUF1_9 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_1_DFFSR_101 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_21_DFFPOSX1_30 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_42_DFFSR_132 INVX1_3/gnd DFFSR_79/S FILL
XFILL_35_DFFSR_63 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_46_DFFSR_23 AND2X2_38/B DFFSR_23/S FILL
XFILL_5_DFFSR_208 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_32_DFFSR_135 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_5_NAND3X1_233 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_46_DFFSR_239 INVX1_39/gnd DFFSR_54/S FILL
XFILL_8_CLKBUF1_3 BUFX2_98/A DFFSR_6/S FILL
XFILL_22_DFFSR_138 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_36_DFFSR_242 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_2_DFFSR_20 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_19_DFFSR_13 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_12_DFFSR_141 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_6_BUFX2_48 AND2X2_38/B DFFSR_59/S FILL
XFILL_26_DFFSR_245 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_16_DFFSR_248 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_1_NOR2X1_1 BUFX2_99/A DFFSR_92/S FILL
XFILL_6_NAND3X1_167 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_43_DFFSR_70 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_8_DFFSR_135 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_49_DFFSR_166 AND2X2_38/B DFFSR_59/S FILL
XNAND3X1_203 NAND3X1_203/A OAI21X1_67/Y OAI21X1_66/Y INVX1_1/gnd AOI22X1_26/D DFFSR_97/S
+ NAND3X1
XFILL_1_INVX1_112 AND2X2_38/B DFFSR_23/S FILL
XFILL_17_CLKBUF1_12 AND2X2_38/B DFFSR_23/S FILL
XFILL_39_DFFSR_169 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_16_DFFSR_60 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_27_DFFSR_20 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_7_NAND3X1_101 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_3_BUFX2_95 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_2_DFFSR_245 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_16_CLKBUF1_15 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_29_DFFSR_172 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_43_DFFSR_276 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_19_DFFSR_175 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_15_CLKBUF1_18 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_33_DFFSR_279 BUFX2_99/A DFFSR_7/S FILL
XFILL_49_1_2 OR2X2_3/gnd DFFSR_4/S FILL
XNOR2X1_57 NOR2X1_57/A NOR2X1_57/B XOR2X1_4/gnd NOR2X1_57/Y DFFSR_91/S NOR2X1
XFILL_14_CLKBUF1_21 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_3_DFFSR_8 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_13_CLKBUF1_24 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_5_XOR2X1_14 INVX1_1/gnd DFFSR_53/S FILL
XFILL_4_NOR2X1_54 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_6_OAI21X1_2 BUFX2_79/A DFFSR_7/S FILL
XFILL_12_CLKBUF1_27 INVX1_1/gnd DFFSR_97/S FILL
XFILL_7_OAI21X1_119 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_35_DFFSR_27 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_7_DFFSR_74 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_11_CLKBUF1_30 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_24_DFFSR_67 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_5_DFFSR_172 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_10_CLKBUF1_33 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_5_NAND3X1_197 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_46_DFFSR_203 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_22_DFFSR_102 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_9_DFFSR_279 BUFX2_99/A DFFSR_7/S FILL
XFILL_1_DFFPOSX1_16 INVX1_67/gnd DFFSR_175/S FILL
XFILL_36_DFFSR_206 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_1_AND2X2_16 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_6_BUFX2_12 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_12_DFFSR_105 INVX1_1/gnd DFFSR_53/S FILL
XFILL_17_0_0 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_26_DFFSR_209 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_9_CLKBUF1_36 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_16_DFFSR_212 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_8_CLKBUF1_39 INVX1_1/gnd DFFSR_53/S FILL
XFILL_6_NAND3X1_131 AND2X2_38/B DFFSR_59/S FILL
XFILL_15_2_1 INVX1_39/gnd DFFSR_34/S FILL
XFILL_7_CLKBUF1_42 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_19_CLKBUF1_7 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_10_DFFPOSX1_35 INVX1_39/gnd DFFSR_54/S FILL
XFILL_4_INVX1_68 INVX1_67/gnd DFFSR_201/S FILL
XFILL_32_DFFSR_74 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_43_DFFSR_34 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_6_CLKBUF1_45 BUFX2_79/A DFFSR_7/S FILL
XFILL_49_DFFSR_130 BUFX2_79/A DFFSR_6/S FILL
XFILL_13_4_2 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_5_CLKBUF1_48 INVX1_3/gnd DFFSR_79/S FILL
XNAND3X1_167 AOI21X1_26/C NAND3X1_167/B INVX1_149/Y XOR2X1_1/gnd NAND2X1_79/B DFFSR_208/S
+ NAND3X1
XFILL_39_DFFSR_133 BUFX2_77/gnd DFFSR_5/S FILL
XCLKBUF1_45 clk BUFX2_79/A CLKBUF1_45/Y DFFSR_7/S CLKBUF1
XFILL_16_DFFSR_24 BUFX2_98/A DFFSR_6/S FILL
XFILL_2_DFFSR_209 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_3_BUFX2_59 AND2X2_38/B DFFSR_23/S FILL
XFILL_29_DFFSR_136 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_43_DFFSR_240 INVX1_39/gnd DFFSR_34/S FILL
XFILL_5_CLKBUF1_4 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_20_DFFPOSX1_24 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_19_DFFSR_139 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_7_NOR3X1_5 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_33_DFFSR_243 BUFX2_7/gnd DFFSR_151/S FILL
XNOR2X1_21 NOR2X1_21/A NOR2X1_21/B DFFSR_28/gnd NOR2X1_21/Y DFFSR_3/S NOR2X1
XFILL_48_DFFSR_8 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_23_DFFSR_246 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_4_NAND3X1_227 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_40_DFFSR_81 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_4_NOR2X1_18 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_13_DFFSR_249 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_0_DFFPOSX1_46 INVX1_39/gnd DFFSR_34/S FILL
XFILL_50_8 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_7_DFFSR_38 BUFX2_98/A DFFSR_6/S FILL
XFILL_24_DFFSR_31 BUFX2_79/A DFFSR_6/S FILL
XFILL_13_DFFSR_71 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_5_DFFSR_136 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_46_DFFSR_167 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_5_NAND3X1_161 AND2X2_38/B DFFSR_23/S FILL
XFILL_9_DFFSR_243 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_36_DFFSR_170 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_50_DFFSR_274 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_0_XOR2X1_8 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_26_DFFSR_173 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_40_DFFSR_277 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_48_DFFSR_88 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_16_DFFSR_176 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_8_AOI22X1_8 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_30_DFFSR_280 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_4_INVX1_32 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_4_DFFSR_85 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_21_DFFSR_78 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_32_DFFSR_38 BUFX2_98/A DFFSR_6/S FILL
XFILL_2_XOR2X1_15 BUFX2_99/A DFFSR_7/S FILL
XFILL_1_NOR2X1_55 INVX1_39/gnd DFFSR_54/S FILL
XFILL_3_OAI21X1_3 BUFX2_99/A DFFSR_92/S FILL
XFILL_5_CLKBUF1_12 AND2X2_38/B DFFSR_23/S FILL
XNAND3X1_131 INVX1_125/Y INVX1_126/Y INVX1_127/Y AND2X2_38/B NAND2X1_55/B DFFSR_59/S
+ NAND3X1
XFILL_4_CLKBUF1_15 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_2_DFFSR_173 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_3_BUFX2_23 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_3_0_2 INVX1_67/gnd DFFSR_175/S FILL
XFILL_29_DFFSR_100 INVX1_1/gnd DFFSR_97/S FILL
XFILL_43_DFFSR_204 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_3_CLKBUF1_18 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_8_AND2X2_14 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_19_DFFSR_103 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_6_DFFSR_280 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_6_OAI21X1_113 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_2_CLKBUF1_21 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_33_DFFSR_207 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_14_DFFSR_6 BUFX2_79/A DFFSR_6/S FILL
XFILL_13_NOR3X1_2 INVX1_1/gnd DFFSR_53/S FILL
XFILL_23_DFFSR_210 BUFX2_98/A DFFSR_6/S FILL
XFILL_4_NAND3X1_191 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_1_CLKBUF1_24 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_40_DFFSR_45 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_1_INVX1_79 INVX1_39/gnd DFFSR_54/S FILL
XFILL_29_DFFSR_85 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_0_DFFPOSX1_10 INVX1_67/gnd DFFSR_201/S FILL
XFILL_0_CLKBUF1_27 INVX1_1/gnd DFFSR_97/S FILL
XFILL_13_DFFSR_213 INVX1_3/gnd DFFSR_23/S FILL
XFILL_16_CLKBUF1_8 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_13_DFFSR_35 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_50_2_0 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_5_DFFSR_100 INVX1_1/gnd DFFSR_97/S FILL
XFILL_0_BUFX2_70 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_5_NAND3X1_125 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_46_DFFSR_131 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_9_DFFSR_207 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_36_DFFSR_134 INVX1_1/gnd DFFSR_53/S FILL
XFILL_48_4_1 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_50_DFFSR_238 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_26_DFFSR_137 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_35_DFFSR_2 BUFX2_79/A DFFSR_7/S FILL
XFILL_10_5 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_40_DFFSR_241 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_2_INVX1_184 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_48_DFFSR_52 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_37_DFFSR_92 BUFX2_99/A DFFSR_92/S FILL
XFILL_2_CLKBUF1_5 BUFX2_99/A DFFSR_92/S FILL
XFILL_16_DFFSR_140 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_46_6_2 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_30_DFFSR_244 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_20_DFFSR_247 BUFX2_99/A DFFSR_7/S FILL
XFILL_10_DFFSR_82 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_21_DFFSR_42 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_4_DFFSR_49 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_19_DFFPOSX1_18 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_1_NOR2X1_19 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_10_DFFSR_250 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_3_NAND3X1_221 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_2_DFFSR_137 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_27_DFFPOSX1_6 AND2X2_38/B DFFSR_23/S FILL
XFILL_43_DFFSR_168 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_45_DFFSR_99 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_26_DFFPOSX1_9 INVX1_67/gnd DFFSR_201/S FILL
XFILL_6_DFFSR_244 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_33_DFFSR_171 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_14_5_0 INVX1_39/gnd DFFSR_54/S FILL
XFILL_47_DFFSR_275 BUFX2_99/A DFFSR_92/S FILL
XFILL_23_DFFSR_174 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_4_NAND3X1_155 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_6_AND2X2_8 BUFX2_99/A DFFSR_7/S FILL
XFILL_1_INVX1_43 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_1_DFFSR_96 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_37_DFFSR_278 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_29_DFFSR_49 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_18_DFFSR_89 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_13_DFFSR_177 DFFSR_46/gnd DFFSR_54/S FILL
XOAI21X1_113 INVX1_211/A NOR2X1_78/Y NAND2X1_173/Y NOR3X1_6/gnd AOI21X1_64/A DFFSR_79/S
+ OAI21X1
XFILL_9_DFFPOSX1_29 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_5_AOI22X1_9 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_9_XOR2X1_13 INVX1_1/gnd DFFSR_97/S FILL
XFILL_0_BUFX2_34 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_0_OAI21X1_4 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_9_DFFSR_171 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_18_DFFPOSX1_48 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_50_DFFSR_202 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_26_DFFSR_101 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_2_INVX1_148 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_40_DFFSR_205 INVX1_3/gnd DFFSR_79/S FILL
XFILL_48_DFFSR_16 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_37_DFFSR_56 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_26_DFFSR_96 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_5_AND2X2_15 INVX1_3/gnd DFFSR_23/S FILL
XFILL_16_DFFSR_104 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_30_DFFSR_208 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_20_DFFSR_211 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_4_DFFSR_13 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_10_DFFSR_46 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_5_OAI21X1_107 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_10_DFFSR_214 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_3_NAND3X1_185 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_13_CLKBUF1_9 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_2_DFFSR_101 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_2_DFFSR_5 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_24_0_0 AND2X2_38/B DFFSR_59/S FILL
XFILL_43_DFFSR_132 INVX1_3/gnd DFFSR_79/S FILL
XFILL_45_DFFSR_63 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_6_DFFSR_208 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_33_DFFSR_135 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_47_DFFSR_239 INVX1_39/gnd DFFSR_54/S FILL
XFILL_9_CLKBUF1_3 BUFX2_98/A DFFSR_6/S FILL
XFILL_22_2_1 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_23_DFFSR_138 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_4_NAND3X1_119 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_37_DFFSR_242 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_1_DFFSR_60 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_29_DFFSR_13 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_18_DFFSR_53 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_4_1_0 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_13_DFFSR_141 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_5_BUFX2_88 INVX1_3/gnd DFFSR_23/S FILL
XFILL_27_DFFSR_245 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_6_NAND2X1_155 BUFX2_79/A DFFSR_7/S FILL
XFILL_0_OR2X2_5 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_20_4_2 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_17_DFFSR_248 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_2_3_1 INVX1_67/gnd DFFSR_201/S FILL
XFILL_26_DFFSR_9 BUFX2_79/A DFFSR_6/S FILL
XFILL_9_DFFSR_135 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_18_DFFPOSX1_12 AND2X2_38/B DFFSR_23/S FILL
XFILL_50_DFFSR_166 AND2X2_38/B DFFSR_59/S FILL
XFILL_0_5_2 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_2_INVX1_112 AND2X2_38/B DFFSR_23/S FILL
XFILL_40_DFFSR_169 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_26_DFFSR_60 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_37_DFFSR_20 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_9_DFFSR_67 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_2_NAND3X1_215 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_3_DFFSR_245 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_30_DFFSR_172 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_44_DFFSR_276 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_20_DFFSR_175 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_10_DFFSR_10 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_34_DFFSR_279 BUFX2_99/A DFFSR_7/S FILL
XFILL_16_DFFPOSX1_3 INVX1_39/gnd DFFSR_34/S FILL
XFILL_10_DFFSR_178 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_15_DFFPOSX1_6 AND2X2_38/B DFFSR_23/S FILL
XFILL_6_XOR2X1_14 INVX1_1/gnd DFFSR_53/S FILL
XFILL_5_NOR2X1_54 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_3_NAND3X1_149 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_47_DFFSR_5 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_14_DFFPOSX1_9 INVX1_67/gnd DFFSR_201/S FILL
XFILL_7_OAI21X1_2 BUFX2_79/A DFFSR_7/S FILL
XFILL_8_DFFPOSX1_23 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_45_DFFSR_27 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_34_DFFSR_67 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_6_DFFSR_172 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_47_DFFSR_203 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_23_DFFSR_102 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_37_DFFSR_206 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_1_DFFSR_24 BUFX2_98/A DFFSR_6/S FILL
XFILL_18_DFFSR_17 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_2_AND2X2_16 NOR3X1_6/gnd DFFSR_91/S FILL
XBUFX2_92 BUFX2_92/A XOR2X1_1/gnd BUFX2_92/Y DFFSR_151/S BUFX2
XFILL_13_DFFSR_105 INVX1_1/gnd DFFSR_53/S FILL
XFILL_5_BUFX2_52 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_27_DFFSR_209 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_17_DFFPOSX1_42 INVX1_39/gnd DFFSR_34/S FILL
XFILL_6_NAND2X1_119 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_2_INVX1_7 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_17_DFFSR_212 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_1_NAND3X1_245 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_0_NOR2X1_5 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_20_CLKBUF1_7 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_9_AOI21X1_44 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_42_DFFSR_74 DFFSR_5/gnd DFFSR_5/S FILL
XNAND2X1_155 DFFSR_7/S NAND2X1_156/A BUFX2_79/A AOI21X1_53/B DFFSR_7/S NAND2X1
XFILL_50_DFFSR_130 BUFX2_79/A DFFSR_6/S FILL
XFILL_4_OAI21X1_101 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_8_AOI21X1_47 INVX1_67/gnd DFFSR_175/S FILL
XFILL_27_DFFPOSX1_31 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_40_DFFSR_133 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_7_AOI21X1_50 INVX1_67/gnd DFFSR_175/S FILL
XFILL_26_DFFSR_24 BUFX2_98/A DFFSR_6/S FILL
XFILL_9_DFFSR_31 BUFX2_79/A DFFSR_6/S FILL
XFILL_15_DFFSR_64 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_2_NAND3X1_179 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_3_DFFSR_209 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_2_BUFX2_99 BUFX2_99/A DFFSR_7/S FILL
XFILL_30_DFFSR_136 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_6_AOI21X1_53 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_44_DFFSR_240 INVX1_39/gnd DFFSR_34/S FILL
XFILL_6_CLKBUF1_4 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_20_DFFSR_139 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_34_DFFSR_243 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_5_AOI21X1_56 NOR3X1_6/gnd DFFSR_79/S FILL
XAOI21X1_53 AOI21X1_53/A AOI21X1_53/B BUFX2_40/Y DFFSR_8/gnd AOI21X1_53/Y DFFSR_60/S
+ AOI21X1
XFILL_10_DFFSR_142 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_4_AOI21X1_59 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_2_XOR2X1_1 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_24_DFFSR_246 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_5_NOR2X1_18 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_13_DFFSR_3 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_50_DFFSR_81 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_3_NAND3X1_113 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_3_AOI21X1_62 INVX1_3/gnd DFFSR_23/S FILL
XFILL_14_DFFSR_249 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_2_AOI21X1_65 INVX1_3/gnd DFFSR_23/S FILL
XFILL_54_5 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_5_NAND2X1_149 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_6_DFFSR_78 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_34_DFFSR_31 BUFX2_79/A DFFSR_6/S FILL
XFILL_23_DFFSR_71 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_6_DFFSR_136 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_1_AOI21X1_68 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_47_DFFSR_167 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_53_6_2 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_0_AOI21X1_71 BUFX2_99/A DFFSR_92/S FILL
XFILL_37_DFFSR_170 OR2X2_6/gnd DFFSR_92/S FILL
XBUFX2_56 BUFX2_58/A BUFX2_8/gnd BUFX2_56/Y DFFSR_51/S BUFX2
XFILL_5_BUFX2_16 BUFX2_98/A DFFSR_32/S FILL
XFILL_0_DFFSR_246 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_27_DFFSR_173 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_41_DFFSR_277 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_17_DFFSR_176 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_8_OAI21X1_95 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_31_DFFSR_280 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_9_AOI22X1_8 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_1_NAND3X1_209 DFFSR_46/gnd DFFSR_62/S FILL
XOAI21X1_6 INVX1_44/Y OAI21X1_4/B OAI21X1_6/C OR2X2_4/gnd NOR2X1_22/B DFFSR_3/S OAI21X1
XFILL_7_OAI21X1_98 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_31_DFFSR_78 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_42_DFFSR_38 BUFX2_98/A DFFSR_6/S FILL
XFILL_3_INVX1_72 NOR3X1_6/gnd DFFSR_79/S FILL
XNAND2X1_119 DFFSR_260/S din[3] DFFSR_5/gnd OAI21X1_88/C DFFSR_5/S NAND2X1
XFILL_3_XOR2X1_15 BUFX2_99/A DFFSR_7/S FILL
XFILL_2_NOR2X1_55 INVX1_39/gnd DFFSR_54/S FILL
XFILL_4_OAI21X1_3 BUFX2_99/A DFFSR_92/S FILL
XFILL_8_AOI21X1_11 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_21_5_0 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_15_DFFSR_28 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_7_AOI21X1_14 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_2_NAND3X1_143 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_3_DFFSR_173 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_2_BUFX2_63 BUFX2_98/A DFFSR_32/S FILL
XFILL_30_DFFSR_100 INVX1_1/gnd DFFSR_97/S FILL
XFILL_6_AOI21X1_17 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_44_DFFSR_204 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_9_AND2X2_14 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_20_DFFSR_103 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_7_DFFSR_280 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_7_DFFPOSX1_17 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_4_DFFPOSX1_3 INVX1_39/gnd DFFSR_34/S FILL
XFILL_4_NAND2X1_179 INVX1_1/gnd DFFSR_97/S FILL
XFILL_5_AOI21X1_20 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_34_DFFSR_207 DFFSR_62/gnd DFFSR_62/S FILL
XAOI21X1_17 INVX1_147/Y NOR3X1_5/A INVX1_148/A BUFX2_7/gnd AOI21X1_17/Y DFFSR_151/S
+ AOI21X1
XFILL_1_6_0 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_10_DFFSR_106 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_3_DFFPOSX1_6 AND2X2_38/B DFFSR_23/S FILL
XFILL_4_AOI21X1_23 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_24_DFFSR_210 BUFX2_98/A DFFSR_6/S FILL
XFILL_50_DFFSR_45 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_39_DFFSR_85 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_2_DFFPOSX1_9 INVX1_67/gnd DFFSR_201/S FILL
XFILL_3_AOI21X1_26 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_14_DFFSR_213 INVX1_3/gnd DFFSR_23/S FILL
XFILL_2_AOI21X1_29 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_16_DFFPOSX1_36 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_17_CLKBUF1_8 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_5_NAND2X1_113 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_6_DFFSR_42 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_23_DFFSR_35 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_6_DFFSR_100 INVX1_1/gnd DFFSR_97/S FILL
XFILL_12_DFFSR_75 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_1_AOI21X1_32 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_0_NAND3X1_239 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_47_DFFSR_131 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_0_AOI21X1_35 INVX1_39/gnd DFFSR_54/S FILL
XFILL_37_DFFSR_134 INVX1_1/gnd DFFSR_53/S FILL
XBUFX2_20 AND2X2_4/Y OR2X2_4/gnd BUFX2_20/Y DFFSR_32/S BUFX2
XFILL_0_DFFSR_210 BUFX2_98/A DFFSR_6/S FILL
XFILL_14_2 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_27_DFFSR_137 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_41_DFFSR_241 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_26_DFFPOSX1_25 BUFX2_79/A DFFSR_6/S FILL
XFILL_3_INVX1_184 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_47_DFFSR_92 BUFX2_99/A DFFSR_92/S FILL
XFILL_3_CLKBUF1_5 BUFX2_99/A DFFSR_92/S FILL
XFILL_17_DFFSR_140 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_31_DFFSR_244 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_8_OAI21X1_59 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_1_NAND3X1_173 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_8_AND2X2_1 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_7_OAI21X1_62 INVX1_3/gnd DFFSR_79/S FILL
XFILL_6_NAND2X1_80 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_21_DFFSR_247 BUFX2_99/A DFFSR_7/S FILL
XFILL_3_INVX1_36 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_31_DFFSR_42 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_31_0_0 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_3_DFFSR_89 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_2_NOR2X1_19 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_20_DFFSR_82 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_6_DFFPOSX1_47 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_6_OAI21X1_65 INVX1_1/gnd DFFSR_53/S FILL
XFILL_5_NAND2X1_83 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_11_DFFSR_250 DFFSR_8/gnd DFFSR_8/S FILL
XNAND2X1_80 INVX1_154/Y NAND2X1_79/Y XOR2X1_1/gnd NAND2X1_80/Y DFFSR_208/S NAND2X1
XFILL_5_OAI21X1_68 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_4_NAND2X1_86 NOR3X1_6/gnd DFFSR_91/S FILL
XOAI21X1_65 INVX1_168/A NOR2X1_71/Y INVX1_167/A INVX1_1/gnd OAI21X1_65/Y DFFSR_53/S
+ OAI21X1
XFILL_29_2_1 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_2_NAND3X1_107 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_3_DFFSR_137 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_4_OAI21X1_71 INVX1_3/gnd DFFSR_79/S FILL
XFILL_3_NAND2X1_89 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_2_BUFX2_27 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_44_DFFSR_168 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_2_NAND2X1_92 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_3_OAI21X1_74 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_1_DFFSR_2 BUFX2_79/A DFFSR_7/S FILL
XFILL_7_DFFSR_244 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_4_NAND2X1_143 INVX1_67/gnd DFFSR_201/S FILL
XFILL_27_4_2 INVX1_3/gnd DFFSR_79/S FILL
XFILL_34_DFFSR_171 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_1_NAND2X1_95 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_12_NOR3X1_6 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_2_OAI21X1_77 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_48_DFFSR_275 BUFX2_99/A DFFSR_92/S FILL
XFILL_24_DFFSR_174 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_1_OAI21X1_80 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_0_NAND2X1_98 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_9_3_1 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_38_DFFSR_278 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_39_DFFSR_49 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_28_DFFSR_89 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_0_INVX1_83 INVX1_39/gnd DFFSR_54/S FILL
XFILL_14_DFFSR_177 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_0_OAI21X1_83 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_6_AOI22X1_9 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_7_5_2 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_12_DFFSR_39 INVX1_3/gnd DFFSR_79/S FILL
XFILL_1_OAI21X1_4 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_0_NAND3X1_203 INVX1_1/gnd DFFSR_97/S FILL
XFILL_51_DFFSR_202 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_0_DFFSR_174 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_27_DFFSR_101 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_25_DFFSR_6 BUFX2_79/A DFFSR_6/S FILL
XFILL_3_INVX1_148 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_41_DFFSR_205 INVX1_3/gnd DFFSR_79/S FILL
XFILL_9_OAI21X1_20 AND2X2_38/B DFFSR_23/S FILL
XFILL_47_DFFSR_56 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_36_DFFSR_96 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_6_AND2X2_15 INVX1_3/gnd DFFSR_23/S FILL
XFILL_17_DFFSR_104 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_8_OAI21X1_23 INVX1_67/gnd DFFSR_201/S FILL
XFILL_31_DFFSR_208 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_1_NAND3X1_137 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_7_OAI21X1_26 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_6_NAND2X1_44 INVX1_39/gnd DFFSR_34/S FILL
XFILL_21_DFFSR_211 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_3_DFFSR_53 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_6_DFFPOSX1_11 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_20_DFFSR_46 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_6_OAI21X1_29 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_5_NAND2X1_47 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_11_DFFSR_214 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_3_NAND2X1_173 NOR3X1_6/gnd DFFSR_79/S FILL
XNAND2X1_44 DFFSR_164/Q AND2X2_18/Y INVX1_39/gnd NAND2X1_44/Y DFFSR_34/S NAND2X1
XFILL_5_OAI21X1_32 AND2X2_38/B DFFSR_59/S FILL
XFILL_4_NAND2X1_50 DFFSR_62/gnd DFFSR_62/S FILL
XOAI21X1_29 INVX1_153/A AND2X2_30/B INVX1_141/A OR2X2_2/gnd XOR2X1_3/B DFFSR_175/S
+ OAI21X1
XFILL_14_CLKBUF1_9 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_4_OAI21X1_35 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_3_DFFSR_101 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_3_NAND2X1_53 DFFSR_62/gnd DFFSR_62/S FILL
XDFFPOSX1_47 AND2X2_33/B CLKBUF1_45/Y AOI21X1_67/Y XOR2X1_4/gnd DFFSR_91/S DFFPOSX1
XFILL_44_DFFSR_132 INVX1_3/gnd DFFSR_79/S FILL
XFILL_15_DFFPOSX1_30 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_2_NAND2X1_56 AND2X2_38/B DFFSR_59/S FILL
XFILL_3_OAI21X1_38 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_46_DFFSR_2 BUFX2_79/A DFFSR_7/S FILL
XFILL_7_DFFSR_208 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_4_NAND2X1_107 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_34_DFFSR_135 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_2_OAI21X1_41 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_1_NAND2X1_59 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_48_DFFSR_239 INVX1_39/gnd DFFSR_54/S FILL
XFILL_24_DFFSR_138 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_38_DFFSR_242 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_0_NAND2X1_62 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_1_OAI21X1_44 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_17_DFFSR_93 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_0_INVX1_185 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_0_INVX1_47 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_39_DFFSR_13 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_28_DFFSR_53 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_10_AOI22X1_10 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_14_DFFSR_141 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_0_CLKBUF1_6 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_19_7 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_0_OAI21X1_47 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_36_2 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_28_DFFSR_245 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_18_DFFSR_248 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_25_DFFPOSX1_19 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_9_AOI22X1_13 AND2X2_38/B DFFSR_23/S FILL
XFILL_0_NAND3X1_167 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_8_AOI22X1_16 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_1_INVX1_4 BUFX2_99/A DFFSR_7/S FILL
XFILL_7_AOI22X1_19 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_5_DFFPOSX1_41 DFFSR_8/gnd DFFSR_60/S FILL
XDFFSR_248 INVX1_117/A DFFSR_3/CLK BUFX2_65/Y DFFSR_8/S DFFSR_240/Q DFFSR_28/gnd DFFSR_8/S
+ DFFSR
XFILL_0_DFFSR_138 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_6_AOI22X1_22 INVX1_3/gnd DFFSR_79/S FILL
XFILL_3_INVX1_112 AND2X2_38/B DFFSR_23/S FILL
XFILL_41_DFFSR_169 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_36_DFFSR_60 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_47_DFFSR_20 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_5_AOI22X1_25 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_4_DFFSR_245 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_31_DFFSR_172 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_1_NAND3X1_101 XOR2X1_4/gnd DFFSR_91/S FILL
XAOI22X1_22 BUFX2_58/Y AND2X2_33/B INVX1_135/A AND2X2_34/B INVX1_3/gnd OAI22X1_50/D
+ DFFSR_79/S AOI22X1
XFILL_45_DFFSR_276 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_4_AOI22X1_28 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_21_DFFSR_175 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_3_DFFSR_17 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_20_DFFSR_10 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_35_DFFSR_279 BUFX2_99/A DFFSR_7/S FILL
XFILL_5_NAND2X1_11 BUFX2_98/A DFFSR_6/S FILL
XFILL_11_DFFSR_178 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_3_NAND2X1_137 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_4_NAND2X1_14 BUFX2_98/A DFFSR_32/S FILL
XFILL_7_XOR2X1_14 INVX1_1/gnd DFFSR_53/S FILL
XFILL_6_NOR2X1_54 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_8_OAI21X1_2 BUFX2_79/A DFFSR_7/S FILL
XFILL_3_NAND2X1_17 OR2X2_6/gnd DFFSR_92/S FILL
XDFFPOSX1_11 OR2X2_1/A CLKBUF1_46/Y NOR2X1_63/Y DFFSR_4/gnd DFFSR_4/S DFFPOSX1
XFILL_2_NAND2X1_20 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_1_OAI21X1_119 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_44_DFFSR_67 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_24_DFFPOSX1_49 BUFX2_99/A DFFSR_92/S FILL
XFILL_7_DFFSR_172 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_1_NAND2X1_23 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_48_DFFSR_203 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_24_DFFSR_102 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_8_NAND3X1_79 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_38_DFFSR_206 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_0_NAND2X1_26 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_0_INVX1_149 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_28_DFFSR_17 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_0_DFFSR_64 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_0_INVX1_11 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_17_DFFSR_57 BUFX2_79/A DFFSR_6/S FILL
XFILL_3_AND2X2_16 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_4_BUFX2_92 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_14_DFFSR_105 INVX1_1/gnd DFFSR_53/S FILL
XFILL_7_NAND3X1_82 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_0_OAI21X1_11 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_28_DFFSR_209 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_6_NAND3X1_85 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_18_DFFSR_212 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_28_5_0 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_5_NAND3X1_88 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_0_NAND3X1_131 AND2X2_38/B DFFSR_59/S FILL
XNAND3X1_85 DFFSR_195/D BUFX2_34/Y BUFX2_23/Y DFFSR_46/gnd NAND3X1_87/A DFFSR_62/S
+ NAND3X1
XFILL_4_NAND3X1_91 AND2X2_38/B DFFSR_59/S FILL
XFILL_3_NAND3X1_94 DFFSR_62/gnd DFFSR_208/S FILL
XDFFSR_212 INVX1_85/A CLKBUF1_31/Y BUFX2_60/Y DFFSR_175/S INVX1_86/A OR2X2_2/gnd DFFSR_175/S
+ DFFSR
XFILL_0_DFFSR_102 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_2_NAND2X1_167 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_8_6_0 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_41_DFFSR_133 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_2_NAND3X1_97 AND2X2_38/B DFFSR_59/S FILL
XFILL_36_DFFSR_24 BUFX2_98/A DFFSR_6/S FILL
XFILL_8_DFFSR_71 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_25_DFFSR_64 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_4_DFFSR_209 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_31_DFFSR_136 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_45_DFFSR_240 INVX1_39/gnd DFFSR_34/S FILL
XFILL_7_CLKBUF1_4 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_21_DFFSR_139 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_35_DFFSR_243 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_14_DFFPOSX1_24 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_11_DFFSR_142 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_3_NAND2X1_101 INVX1_39/gnd DFFSR_54/S FILL
XFILL_25_DFFSR_246 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_6_NOR2X1_18 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_15_DFFSR_249 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_37_DFFSR_9 BUFX2_79/A DFFSR_6/S FILL
XFILL_11_OAI22X1_19 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_10_OAI22X1_22 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_44_DFFSR_31 BUFX2_79/A DFFSR_6/S FILL
XFILL_33_DFFSR_71 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_7_DFFSR_136 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_24_DFFPOSX1_13 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_48_DFFSR_167 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_8_NAND3X1_43 BUFX2_99/A DFFSR_7/S FILL
XFILL_9_OAI22X1_25 INVX1_39/gnd DFFSR_54/S FILL
XFILL_38_DFFSR_170 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_0_DFFSR_28 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_0_INVX1_113 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_17_DFFSR_21 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_8_NAND3X1_216 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_7_NAND3X1_46 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_38_0_0 BUFX2_79/A DFFSR_7/S FILL
XFILL_8_OAI22X1_28 INVX1_3/gnd DFFSR_23/S FILL
XFILL_4_BUFX2_56 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_1_DFFSR_246 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_28_DFFSR_173 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_4_DFFPOSX1_35 INVX1_39/gnd DFFSR_54/S FILL
XFILL_42_DFFSR_277 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_6_NAND3X1_49 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_7_OAI22X1_31 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_18_DFFSR_176 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_8_NOR3X1_2 INVX1_1/gnd DFFSR_53/S FILL
XFILL_5_NAND3X1_52 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_32_DFFSR_280 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_36_2_1 BUFX2_99/A DFFSR_92/S FILL
XFILL_6_OAI22X1_34 DFFSR_34/gnd DFFSR_1/S FILL
XNAND3X1_49 DFFSR_63/D BUFX2_17/Y BUFX2_13/Y DFFSR_8/gnd NAND3X1_49/Y DFFSR_60/S NAND3X1
XFILL_4_NAND3X1_55 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_5_OAI22X1_37 INVX1_3/gnd DFFSR_23/S FILL
XFILL_41_DFFSR_78 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_4_XOR2X1_15 BUFX2_99/A DFFSR_7/S FILL
XFILL_3_NOR2X1_55 INVX1_39/gnd DFFSR_54/S FILL
XOAI22X1_34 INVX1_83/Y OAI22X1_43/B INVX1_84/Y OAI22X1_43/D DFFSR_34/gnd NOR2X1_44/B
+ DFFSR_1/S OAI22X1
XFILL_3_NAND3X1_58 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_5_OAI21X1_3 BUFX2_99/A DFFSR_92/S FILL
XFILL_4_OAI22X1_40 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_34_4_2 OR2X2_6/gnd DFFSR_53/S FILL
XDFFSR_176 DFFSR_192/D CLKBUF1_39/Y BUFX2_63/Y DFFSR_53/S DFFSR_176/D OR2X2_6/gnd
+ DFFSR_53/S DFFSR
XFILL_2_NAND2X1_131 INVX1_3/gnd DFFSR_79/S FILL
XFILL_2_NAND3X1_61 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_3_OAI22X1_43 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_8_DFFSR_35 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_25_DFFSR_28 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_14_DFFSR_68 BUFX2_98/A DFFSR_6/S FILL
XFILL_4_DFFSR_173 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_31_DFFSR_100 INVX1_1/gnd DFFSR_97/S FILL
XFILL_1_NAND3X1_64 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_2_OAI22X1_46 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_45_DFFSR_204 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_21_DFFSR_103 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_0_NAND3X1_67 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_8_DFFSR_280 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_1_OAI22X1_49 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_35_DFFSR_207 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_0_OAI21X1_113 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_23_DFFPOSX1_43 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_0_AND2X2_17 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_0_OAI22X1_52 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_11_DFFSR_106 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_25_DFFSR_210 BUFX2_98/A DFFSR_6/S FILL
XFILL_1_XOR2X1_5 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_49_DFFSR_85 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_7_NAND3X1_246 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_15_DFFSR_213 INVX1_3/gnd DFFSR_23/S FILL
XFILL_18_CLKBUF1_8 NOR3X1_6/gnd DFFSR_79/S FILL
XINVX1_69 INVX1_69/A INVX1_3/gnd INVX1_69/Y DFFSR_23/S INVX1
XFILL_33_DFFSR_35 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_5_DFFSR_82 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_22_DFFSR_75 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_7_DFFSR_100 INVX1_1/gnd DFFSR_97/S FILL
XFILL_48_DFFSR_131 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_38_DFFSR_134 INVX1_1/gnd DFFSR_53/S FILL
XFILL_8_NAND3X1_180 OR2X2_1/gnd DFFSR_59/S FILL
XINVX1_187 DFFSR_7/D OR2X2_1/gnd INVX1_187/Y DFFSR_59/S INVX1
XFILL_4_BUFX2_20 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_1_DFFSR_210 BUFX2_98/A DFFSR_6/S FILL
XFILL_7_NAND3X1_10 BUFX2_79/A DFFSR_6/S FILL
XCLKBUF1_8 BUFX2_4/Y NOR3X1_6/gnd CLKBUF1_8/Y DFFSR_79/S CLKBUF1
XFILL_28_DFFSR_137 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_42_DFFSR_241 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_1_NAND2X1_161 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_6_NAND3X1_13 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_4_INVX1_184 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_4_CLKBUF1_5 BUFX2_99/A DFFSR_92/S FILL
XFILL_18_DFFSR_140 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_5_NAND3X1_16 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_24_DFFSR_3 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_32_DFFSR_244 DFFSR_1/gnd DFFSR_81/S FILL
XNAND3X1_13 DFFSR_66/D BUFX2_19/Y BUFX2_13/Y DFFSR_4/gnd NAND3X1_13/Y DFFSR_4/S NAND3X1
XFILL_22_DFFSR_247 BUFX2_99/A DFFSR_7/S FILL
XFILL_41_DFFSR_42 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_4_NAND3X1_19 BUFX2_99/A DFFSR_92/S FILL
XFILL_2_INVX1_76 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_30_DFFSR_82 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_3_NOR2X1_19 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_12_DFFSR_250 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_13_DFFPOSX1_18 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_3_NAND3X1_22 OR2X2_6/gnd DFFSR_53/S FILL
XDFFSR_140 DFFSR_196/D CLKBUF1_11/Y BUFX2_68/Y DFFSR_208/S INVX1_83/A DFFSR_62/gnd
+ DFFSR_208/S DFFSR
XFILL_2_NAND3X1_25 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_14_DFFSR_32 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_4_DFFSR_137 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_1_BUFX2_67 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_1_NAND3X1_28 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_2_OAI22X1_10 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_45_DFFSR_168 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_0_NAND3X1_31 BUFX2_79/A DFFSR_6/S FILL
XFILL_1_OAI22X1_13 INVX1_1/gnd DFFSR_53/S FILL
XFILL_8_DFFSR_244 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_35_DFFSR_171 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_49_DFFSR_275 BUFX2_99/A DFFSR_92/S FILL
XFILL_0_OAI22X1_16 AND2X2_38/B DFFSR_59/S FILL
XFILL_25_DFFSR_174 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_49_DFFSR_49 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_38_DFFSR_89 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_39_DFFSR_278 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_7_NAND3X1_210 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_15_DFFSR_177 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_7_AOI22X1_9 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_3_DFFPOSX1_29 BUFX2_72/gnd DFFSR_276/S FILL
XINVX1_33 INVX1_33/A DFFSR_28/gnd INVX1_33/Y DFFSR_3/S INVX1
XDFFSR_86 DFFSR_86/Q DFFSR_45/CLK DFFSR_15/R DFFSR_4/S DFFSR_78/Q DFFSR_4/gnd DFFSR_4/S
+ DFFSR
XFILL_10_0_1 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_22_DFFSR_39 INVX1_3/gnd DFFSR_79/S FILL
XFILL_5_DFFSR_46 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_11_DFFSR_79 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_0_NOR2X1_56 AND2X2_38/B DFFSR_59/S FILL
XFILL_2_OAI21X1_4 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_8_NAND3X1_144 AND2X2_38/B DFFSR_59/S FILL
XINVX1_151 INVX1_151/A OR2X2_1/gnd INVX1_151/Y DFFSR_51/S INVX1
XFILL_0_INVX1_1 INVX1_1/gnd DFFSR_53/S FILL
XFILL_1_3 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_12_DFFPOSX1_48 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_1_DFFSR_174 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_28_DFFSR_101 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_1_NAND2X1_125 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_15_XOR2X1_9 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_42_DFFSR_205 INVX1_3/gnd DFFSR_79/S FILL
XFILL_46_DFFSR_96 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_7_AND2X2_15 INVX1_3/gnd DFFSR_23/S FILL
XFILL_18_DFFSR_104 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_32_DFFSR_208 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_22_DFFSR_211 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_7_AND2X2_5 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_2_INVX1_40 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_2_DFFSR_93 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_19_DFFSR_86 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_30_DFFSR_46 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_12_DFFSR_214 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_22_DFFPOSX1_37 BUFX2_72/gnd DFFSR_201/S FILL
XDFFSR_104 DFFSR_112/D CLKBUF1_7/Y DFFSR_35/R DFFSR_8/S DFFSR_96/Q DFFSR_28/gnd DFFSR_8/S
+ DFFSR
XFILL_15_CLKBUF1_9 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_4_DFFSR_101 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_6_NAND3X1_240 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_1_BUFX2_31 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_45_DFFSR_132 INVX1_3/gnd DFFSR_79/S FILL
XFILL_8_DFFSR_208 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_35_DFFSR_135 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_35_5_0 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_49_DFFSR_239 INVX1_39/gnd DFFSR_54/S FILL
XFILL_25_DFFSR_138 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_39_DFFSR_242 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_1_INVX1_185 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_49_DFFSR_13 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_38_DFFSR_53 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_27_DFFSR_93 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_15_DFFSR_141 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_7_NAND3X1_174 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_1_CLKBUF1_6 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_29_DFFSR_245 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_19_DFFSR_248 DFFSR_28/gnd DFFSR_8/S FILL
XDFFSR_50 DFFSR_50/Q CLKBUF1_37/Y DFFSR_8/R DFFSR_5/S DFFSR_58/Q BUFX2_77/gnd DFFSR_5/S
+ DFFSR
XFILL_0_NAND2X1_155 BUFX2_79/A DFFSR_7/S FILL
XFILL_5_DFFSR_10 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_11_DFFSR_43 BUFX2_98/A DFFSR_6/S FILL
XFILL_0_NOR2X1_20 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_8_NAND3X1_108 BUFX2_8/gnd DFFSR_81/S FILL
XINVX1_115 INVX1_115/A XOR2X1_4/gnd INVX1_115/Y DFFSR_91/S INVX1
XFILL_12_DFFPOSX1_12 AND2X2_38/B DFFSR_23/S FILL
XFILL_1_DFFSR_138 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_42_DFFSR_169 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_4_INVX1_112 AND2X2_38/B DFFSR_23/S FILL
XFILL_46_DFFSR_60 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_5_DFFSR_245 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_32_DFFSR_172 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_46_DFFSR_276 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_22_DFFSR_175 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_2_DFFSR_57 BUFX2_79/A DFFSR_6/S FILL
XFILL_30_DFFSR_10 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_19_DFFSR_50 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_36_DFFSR_279 BUFX2_99/A DFFSR_7/S FILL
XFILL_6_BUFX2_85 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_12_DFFSR_178 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_8_XOR2X1_14 INVX1_1/gnd DFFSR_53/S FILL
XFILL_9_OAI21X1_2 BUFX2_79/A DFFSR_7/S FILL
XFILL_20_CLKBUF1_40 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_6_NAND3X1_204 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_45_0_0 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_36_DFFSR_6 BUFX2_79/A DFFSR_6/S FILL
XFILL_2_DFFPOSX1_23 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_19_CLKBUF1_43 AND2X2_38/B DFFSR_23/S FILL
XFILL_8_DFFSR_172 DFFSR_46/gnd DFFSR_62/S FILL
XAND2X2_19 AND2X2_19/A AND2X2_19/B BUFX2_7/gnd AND2X2_19/Y DFFSR_216/S AND2X2
XFILL_18_CLKBUF1_46 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_49_DFFSR_203 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_25_DFFSR_102 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_43_2_1 OR2X2_4/gnd DFFSR_3/S FILL
XNAND3X1_240 INVX1_179/A NAND3X1_239/A NAND3X1_239/B DFFSR_8/gnd AOI21X1_39/B DFFSR_60/S
+ NAND3X1
XFILL_39_DFFSR_206 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_17_CLKBUF1_49 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_1_INVX1_149 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_38_DFFSR_17 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_27_DFFSR_57 BUFX2_79/A DFFSR_6/S FILL
XFILL_16_DFFSR_97 INVX1_1/gnd DFFSR_97/S FILL
XFILL_4_AND2X2_16 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_7_NAND3X1_138 INVX1_67/gnd DFFSR_201/S FILL
XFILL_15_DFFSR_105 INVX1_1/gnd DFFSR_53/S FILL
XFILL_29_DFFSR_209 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_11_DFFPOSX1_42 INVX1_39/gnd DFFSR_34/S FILL
XFILL_41_4_2 BUFX2_98/A DFFSR_32/S FILL
XFILL_19_DFFSR_212 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_0_NAND2X1_119 DFFSR_5/gnd DFFSR_5/S FILL
XDFFSR_14 DFFSR_14/Q DFFSR_83/CLK DFFSR_7/R DFFSR_53/S DFFSR_54/Q INVX1_1/gnd DFFSR_53/S
+ DFFSR
XFILL_1_DFFSR_102 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_42_DFFSR_133 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_21_DFFPOSX1_31 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_35_DFFSR_64 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_46_DFFSR_24 BUFX2_98/A DFFSR_6/S FILL
XFILL_5_DFFSR_209 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_32_DFFSR_136 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_46_DFFSR_240 INVX1_39/gnd DFFSR_34/S FILL
XFILL_5_NAND3X1_234 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_8_CLKBUF1_4 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_22_DFFSR_139 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_2_DFFSR_21 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_36_DFFSR_243 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_19_DFFSR_14 INVX1_1/gnd DFFSR_53/S FILL
XFILL_12_DFFSR_142 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_6_BUFX2_49 INVX1_1/gnd DFFSR_97/S FILL
XFILL_26_DFFSR_246 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_16_DFFSR_249 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_1_NOR2X1_2 INVX1_1/gnd DFFSR_97/S FILL
XFILL_6_NAND3X1_168 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_43_DFFSR_71 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_8_DFFSR_136 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_18_CLKBUF1_10 INVX1_67/gnd DFFSR_201/S FILL
XFILL_49_DFFSR_167 OR2X2_2/gnd DFFSR_216/S FILL
XNAND3X1_204 NAND3X1_201/A OAI21X1_65/Y OAI21X1_66/Y OR2X2_6/gnd INVX1_174/A DFFSR_53/S
+ NAND3X1
XFILL_17_CLKBUF1_13 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_39_DFFSR_170 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_1_INVX1_113 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_27_DFFSR_21 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_16_DFFSR_61 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_7_NAND3X1_102 INVX1_3/gnd DFFSR_23/S FILL
XFILL_2_DFFSR_246 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_3_BUFX2_96 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_16_CLKBUF1_16 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_29_DFFSR_173 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_43_DFFSR_277 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_19_DFFSR_176 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_15_CLKBUF1_19 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_33_DFFSR_280 OR2X2_6/gnd DFFSR_53/S FILL
XNOR2X1_58 NOR2X1_58/A NOR2X1_58/B INVX1_3/gnd NOR2X1_58/Y DFFSR_79/S NOR2X1
XFILL_14_CLKBUF1_22 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_3_DFFSR_9 BUFX2_79/A DFFSR_6/S FILL
XFILL_51_DFFSR_78 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_5_XOR2X1_15 BUFX2_99/A DFFSR_7/S FILL
XFILL_13_CLKBUF1_25 INVX1_67/gnd DFFSR_201/S FILL
XFILL_4_NOR2X1_55 INVX1_39/gnd DFFSR_54/S FILL
XFILL_6_OAI21X1_3 BUFX2_99/A DFFSR_92/S FILL
XFILL_12_CLKBUF1_28 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_11_CLKBUF1_31 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_35_DFFSR_28 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_24_DFFSR_68 BUFX2_98/A DFFSR_6/S FILL
XFILL_7_DFFSR_75 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_5_DFFSR_173 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_32_DFFSR_100 INVX1_1/gnd DFFSR_97/S FILL
XFILL_10_CLKBUF1_34 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_46_DFFSR_204 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_5_NAND3X1_198 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_22_DFFSR_103 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_9_DFFSR_280 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_1_DFFPOSX1_17 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_36_DFFSR_207 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_1_AND2X2_17 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_17_0_1 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_6_BUFX2_13 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_12_DFFSR_106 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_9_CLKBUF1_37 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_26_DFFSR_210 BUFX2_98/A DFFSR_6/S FILL
XFILL_16_DFFSR_213 INVX1_3/gnd DFFSR_23/S FILL
XFILL_8_CLKBUF1_40 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_6_NAND3X1_132 AND2X2_38/B DFFSR_23/S FILL
XFILL_15_2_2 INVX1_39/gnd DFFSR_34/S FILL
XFILL_7_CLKBUF1_43 AND2X2_38/B DFFSR_23/S FILL
XFILL_10_DFFPOSX1_36 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_19_CLKBUF1_8 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_43_DFFSR_35 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_4_INVX1_69 INVX1_3/gnd DFFSR_23/S FILL
XFILL_8_DFFSR_100 INVX1_1/gnd DFFSR_97/S FILL
XFILL_32_DFFSR_75 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_6_CLKBUF1_46 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_49_DFFSR_131 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_5_CLKBUF1_49 BUFX2_8/gnd DFFSR_81/S FILL
XNAND3X1_168 INVX1_154/A OAI21X1_42/Y NAND2X1_79/B XOR2X1_1/gnd INVX1_156/A DFFSR_208/S
+ NAND3X1
XFILL_39_DFFSR_134 INVX1_1/gnd DFFSR_53/S FILL
XCLKBUF1_46 clk OR2X2_3/gnd CLKBUF1_46/Y DFFSR_4/S CLKBUF1
XFILL_16_DFFSR_25 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_2_DFFSR_210 BUFX2_98/A DFFSR_6/S FILL
XFILL_3_BUFX2_60 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_29_DFFSR_137 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_43_DFFSR_241 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_20_DFFPOSX1_25 BUFX2_79/A DFFSR_6/S FILL
XFILL_5_CLKBUF1_5 BUFX2_99/A DFFSR_92/S FILL
XFILL_19_DFFSR_140 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_7_NOR3X1_6 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_33_DFFSR_244 DFFSR_1/gnd DFFSR_81/S FILL
XNOR2X1_22 NOR2X1_22/A NOR2X1_22/B OR2X2_4/gnd NOR2X1_22/Y DFFSR_3/S NOR2X1
XFILL_48_DFFSR_9 BUFX2_79/A DFFSR_6/S FILL
XFILL_4_NAND3X1_228 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_23_DFFSR_247 BUFX2_99/A DFFSR_7/S FILL
XFILL_40_DFFSR_82 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_51_DFFSR_42 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_4_NOR2X1_19 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_13_DFFSR_250 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_0_DFFPOSX1_47 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_42_5_0 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_50_9 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_13_DFFSR_72 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_24_DFFSR_32 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_7_DFFSR_39 INVX1_3/gnd DFFSR_79/S FILL
XFILL_5_DFFSR_137 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_46_DFFSR_168 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_5_NAND3X1_162 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_9_DFFSR_244 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_36_DFFSR_171 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_50_DFFSR_275 BUFX2_99/A DFFSR_92/S FILL
XFILL_0_XOR2X1_9 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_26_DFFSR_174 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_48_DFFSR_89 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_40_DFFSR_278 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_16_DFFSR_177 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_8_AOI22X1_9 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_4_INVX1_33 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_4_DFFSR_86 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_32_DFFSR_39 INVX1_3/gnd DFFSR_79/S FILL
XFILL_21_DFFSR_79 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_6_CLKBUF1_10 INVX1_67/gnd DFFSR_201/S FILL
XFILL_1_NOR2X1_56 AND2X2_38/B DFFSR_59/S FILL
XFILL_3_OAI21X1_4 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_5_CLKBUF1_13 DFFSR_28/gnd DFFSR_3/S FILL
XNAND3X1_132 INVX1_124/Y OAI21X1_20/Y NAND2X1_55/B AND2X2_38/B DFFPOSX1_8/D DFFSR_23/S
+ NAND3X1
XCLKBUF1_10 BUFX2_5/Y INVX1_67/gnd CLKBUF1_10/Y DFFSR_201/S CLKBUF1
XFILL_4_CLKBUF1_16 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_2_DFFSR_174 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_3_BUFX2_24 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_29_DFFSR_101 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_43_DFFSR_205 INVX1_3/gnd DFFSR_79/S FILL
XFILL_3_CLKBUF1_19 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_8_AND2X2_15 INVX1_3/gnd DFFSR_23/S FILL
XFILL_19_DFFSR_104 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_6_OAI21X1_114 AND2X2_38/B DFFSR_59/S FILL
XFILL_13_NOR3X1_3 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_14_DFFSR_7 BUFX2_79/A DFFSR_7/S FILL
XFILL_2_CLKBUF1_22 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_33_DFFSR_208 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_1_CLKBUF1_25 INVX1_67/gnd DFFSR_201/S FILL
XFILL_4_NAND3X1_192 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_23_DFFSR_211 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_29_DFFSR_86 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_52_0_0 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_1_INVX1_80 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_40_DFFSR_46 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_13_DFFSR_214 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_0_DFFPOSX1_11 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_0_CLKBUF1_28 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_16_CLKBUF1_9 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_50_2_1 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_13_DFFSR_36 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_5_DFFSR_101 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_0_BUFX2_71 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_46_DFFSR_132 INVX1_3/gnd DFFSR_79/S FILL
XFILL_5_NAND3X1_126 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_9_DFFSR_208 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_36_DFFSR_135 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_48_4_2 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_50_DFFSR_239 INVX1_39/gnd DFFSR_54/S FILL
XFILL_35_DFFSR_3 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_26_DFFSR_138 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_10_6 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_40_DFFSR_242 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_2_INVX1_185 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_48_DFFSR_53 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_27_1 INVX1_3/gnd DFFSR_23/S FILL
XFILL_37_DFFSR_93 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_16_DFFSR_141 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_2_CLKBUF1_6 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_30_DFFSR_245 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_20_DFFSR_248 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_4_DFFSR_50 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_21_DFFSR_43 BUFX2_98/A DFFSR_6/S FILL
XFILL_10_DFFSR_83 INVX1_3/gnd DFFSR_79/S FILL
XFILL_19_DFFPOSX1_19 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_1_NOR2X1_20 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_10_DFFSR_251 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_3_NAND3X1_222 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_2_DFFSR_138 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_16_3_0 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_27_DFFPOSX1_7 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_43_DFFSR_169 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_6_DFFSR_245 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_33_DFFSR_172 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_14_5_1 INVX1_39/gnd DFFSR_54/S FILL
XFILL_47_DFFSR_276 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_23_DFFSR_175 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_6_AND2X2_9 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_4_NAND3X1_156 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_40_DFFSR_10 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_29_DFFSR_50 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_1_INVX1_44 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_37_DFFSR_279 BUFX2_99/A DFFSR_7/S FILL
XFILL_1_DFFSR_97 INVX1_1/gnd DFFSR_97/S FILL
XFILL_18_DFFSR_90 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_13_DFFSR_178 NOR3X1_6/gnd DFFSR_79/S FILL
XOAI21X1_114 XOR2X1_10/Y AOI21X1_64/A INVX1_212/Y AND2X2_38/B AOI21X1_64/C DFFSR_59/S
+ OAI21X1
XFILL_9_DFFPOSX1_30 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_9_XOR2X1_14 INVX1_1/gnd DFFSR_53/S FILL
XFILL_0_BUFX2_35 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_0_OAI21X1_5 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_9_DFFSR_172 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_18_DFFPOSX1_49 BUFX2_99/A DFFSR_92/S FILL
XFILL_50_DFFSR_203 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_26_DFFSR_102 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_40_DFFSR_206 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_2_INVX1_149 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_48_DFFSR_17 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_37_DFFSR_57 BUFX2_79/A DFFSR_6/S FILL
XFILL_26_DFFSR_97 INVX1_1/gnd DFFSR_97/S FILL
XFILL_5_AND2X2_16 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_16_DFFSR_105 INVX1_1/gnd DFFSR_53/S FILL
XFILL_30_DFFSR_209 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_20_DFFSR_212 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_4_DFFSR_14 INVX1_1/gnd DFFSR_53/S FILL
XFILL_10_DFFSR_47 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_5_OAI21X1_108 INVX1_1/gnd DFFSR_53/S FILL
XFILL_10_DFFSR_215 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_3_NAND3X1_186 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_2_DFFSR_102 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_2_DFFSR_6 BUFX2_79/A DFFSR_6/S FILL
XFILL_24_0_1 AND2X2_38/B DFFSR_59/S FILL
XFILL_43_DFFSR_133 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_45_DFFSR_64 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_6_DFFSR_209 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_33_DFFSR_136 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_47_DFFSR_240 INVX1_39/gnd DFFSR_34/S FILL
XFILL_9_CLKBUF1_4 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_22_2_2 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_4_NAND3X1_120 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_23_DFFSR_139 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_37_DFFSR_243 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_1_DFFSR_61 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_29_DFFSR_14 INVX1_1/gnd DFFSR_53/S FILL
XFILL_18_DFFSR_54 INVX1_39/gnd DFFSR_54/S FILL
XFILL_13_DFFSR_142 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_4_1_1 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_5_BUFX2_89 INVX1_1/gnd DFFSR_97/S FILL
XFILL_27_DFFSR_246 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_0_OR2X2_6 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_6_NAND2X1_156 AND2X2_38/B DFFSR_59/S FILL
XFILL_17_DFFSR_249 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_49_1 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_2_3_2 INVX1_67/gnd DFFSR_201/S FILL
XFILL_9_DFFSR_136 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_50_DFFSR_167 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_18_DFFPOSX1_13 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_2_INVX1_113 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_9_DFFSR_68 BUFX2_98/A DFFSR_6/S FILL
XFILL_40_DFFSR_170 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_26_DFFSR_61 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_37_DFFSR_21 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_2_NAND3X1_216 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_3_DFFSR_246 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_30_DFFSR_173 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_44_DFFSR_277 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_17_DFFPOSX1_1 INVX1_39/gnd DFFSR_34/S FILL
XFILL_20_DFFSR_176 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_49_5_0 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_34_DFFSR_280 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_10_DFFSR_11 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_16_DFFPOSX1_4 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_10_DFFSR_179 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_15_DFFPOSX1_7 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_6_XOR2X1_15 BUFX2_99/A DFFSR_7/S FILL
XFILL_3_NAND3X1_150 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_5_NOR2X1_55 INVX1_39/gnd DFFSR_54/S FILL
XFILL_47_DFFSR_6 BUFX2_79/A DFFSR_6/S FILL
XFILL_7_OAI21X1_3 BUFX2_99/A DFFSR_92/S FILL
XFILL_8_DFFPOSX1_24 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_45_DFFSR_28 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_34_DFFSR_68 BUFX2_98/A DFFSR_6/S FILL
XFILL_6_DFFSR_173 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_33_DFFSR_100 INVX1_1/gnd DFFSR_97/S FILL
XFILL_47_DFFSR_204 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_23_DFFSR_103 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_1_DFFSR_25 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_18_DFFSR_18 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_37_DFFSR_207 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_2_AND2X2_17 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_13_DFFSR_106 XOR2X1_4/gnd DFFSR_91/S FILL
XBUFX2_93 BUFX2_93/A AND2X2_38/B BUFX2_93/Y DFFSR_59/S BUFX2
XFILL_17_DFFPOSX1_43 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_5_BUFX2_53 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_27_DFFSR_210 BUFX2_98/A DFFSR_6/S FILL
XFILL_6_NAND2X1_120 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_2_INVX1_8 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_17_DFFSR_213 INVX1_3/gnd DFFSR_23/S FILL
XFILL_1_NAND3X1_246 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_0_NOR2X1_6 BUFX2_98/A DFFSR_6/S FILL
XFILL_20_CLKBUF1_8 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_9_DFFSR_100 INVX1_1/gnd DFFSR_97/S FILL
XFILL_42_DFFSR_75 DFFSR_34/gnd DFFSR_1/S FILL
XNAND2X1_156 NAND2X1_156/A INVX1_208/Y AND2X2_38/B AOI21X1_54/A DFFSR_59/S NAND2X1
XFILL_50_DFFSR_131 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_4_OAI21X1_102 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_8_AOI21X1_48 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_27_DFFPOSX1_32 INVX1_67/gnd DFFSR_201/S FILL
XFILL_40_DFFSR_134 INVX1_1/gnd DFFSR_53/S FILL
XFILL_9_DFFSR_32 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_26_DFFSR_25 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_15_DFFSR_65 BUFX2_79/A DFFSR_7/S FILL
XFILL_7_AOI21X1_51 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_3_DFFSR_210 BUFX2_98/A DFFSR_6/S FILL
XFILL_2_NAND3X1_180 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_30_DFFSR_137 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_6_AOI21X1_54 AND2X2_38/B DFFSR_59/S FILL
XFILL_44_DFFSR_241 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_6_CLKBUF1_5 BUFX2_99/A DFFSR_92/S FILL
XFILL_20_DFFSR_140 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_5_AOI21X1_57 INVX1_67/gnd DFFSR_201/S FILL
XFILL_34_DFFSR_244 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_10_DFFSR_143 OR2X2_2/gnd DFFSR_216/S FILL
XAOI21X1_54 AOI21X1_54/A AOI21X1_54/B BUFX2_35/Y AND2X2_38/B AOI21X1_54/Y DFFSR_59/S
+ AOI21X1
XFILL_4_AOI21X1_60 BUFX2_79/A DFFSR_7/S FILL
XFILL_2_XOR2X1_2 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_24_DFFSR_247 BUFX2_99/A DFFSR_7/S FILL
XFILL_50_DFFSR_82 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_5_NOR2X1_19 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_13_DFFSR_4 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_3_NAND3X1_114 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_14_DFFSR_250 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_3_AOI21X1_63 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_2_AOI21X1_66 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_54_6 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_34_DFFSR_32 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_6_DFFSR_79 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_5_NAND2X1_150 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_6_DFFSR_137 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_23_DFFSR_72 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_1_AOI21X1_69 INVX1_1/gnd DFFSR_97/S FILL
XFILL_47_DFFSR_168 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_37_DFFSR_171 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_0_DFFSR_247 BUFX2_99/A DFFSR_7/S FILL
XFILL_51_DFFSR_275 BUFX2_99/A DFFSR_92/S FILL
XBUFX2_57 BUFX2_58/A AND2X2_38/B BUFX2_57/Y DFFSR_23/S BUFX2
XFILL_5_BUFX2_17 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_27_DFFSR_174 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_9_OAI21X1_93 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_41_DFFSR_278 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_17_DFFSR_177 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_9_AOI22X1_9 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_8_OAI21X1_96 AND2X2_38/B DFFSR_59/S FILL
XFILL_1_NAND3X1_210 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_23_3_0 OR2X2_1/gnd DFFSR_59/S FILL
XOAI21X1_7 INVX1_51/Y OAI21X1_4/B OAI21X1_7/C DFFSR_8/gnd NOR2X1_25/B DFFSR_8/S OAI21X1
XFILL_7_OAI21X1_99 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_31_DFFSR_79 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_42_DFFSR_39 INVX1_3/gnd DFFSR_79/S FILL
XFILL_3_INVX1_73 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_2_NOR2X1_56 AND2X2_38/B DFFSR_59/S FILL
XNAND2X1_120 DFFSR_54/S din[4] DFFSR_46/gnd OAI21X1_89/C DFFSR_54/S NAND2X1
XFILL_4_OAI21X1_4 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_8_AOI21X1_12 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_21_5_1 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_15_DFFSR_29 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_7_AOI21X1_15 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_2_NAND3X1_144 AND2X2_38/B DFFSR_59/S FILL
XFILL_3_DFFSR_174 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_3_4_0 INVX1_67/gnd DFFSR_175/S FILL
XFILL_2_BUFX2_64 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_30_DFFSR_101 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_6_AOI21X1_18 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_5_DFFPOSX1_1 INVX1_39/gnd DFFSR_34/S FILL
XFILL_44_DFFSR_205 INVX1_3/gnd DFFSR_79/S FILL
XFILL_9_AND2X2_15 INVX1_3/gnd DFFSR_23/S FILL
XFILL_20_DFFSR_104 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_7_DFFPOSX1_18 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_5_AOI21X1_21 INVX1_39/gnd DFFSR_54/S FILL
XFILL_4_DFFPOSX1_4 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_4_NAND2X1_180 INVX1_1/gnd DFFSR_97/S FILL
XFILL_34_DFFSR_208 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_1_6_1 BUFX2_72/gnd DFFSR_201/S FILL
XAOI21X1_18 AOI21X1_18/A XOR2X1_3/B INVX1_155/Y OR2X2_2/gnd AOI21X1_18/Y DFFSR_175/S
+ AOI21X1
XFILL_10_DFFSR_107 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_3_DFFPOSX1_7 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_4_AOI21X1_24 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_24_DFFSR_211 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_39_DFFSR_86 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_50_DFFSR_46 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_14_DFFSR_214 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_3_AOI21X1_27 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_16_DFFPOSX1_37 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_2_AOI21X1_30 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_17_CLKBUF1_9 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_5_NAND2X1_114 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_6_DFFSR_43 BUFX2_98/A DFFSR_6/S FILL
XFILL_6_DFFSR_101 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_23_DFFSR_36 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_12_DFFSR_76 BUFX2_79/A DFFSR_7/S FILL
XFILL_1_AOI21X1_33 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_0_NAND3X1_240 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_47_DFFSR_132 INVX1_3/gnd DFFSR_79/S FILL
XFILL_0_AOI21X1_36 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_37_DFFSR_135 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_0_DFFSR_211 BUFX2_7/gnd DFFSR_216/S FILL
XBUFX2_21 AND2X2_4/Y OR2X2_4/gnd BUFX2_21/Y DFFSR_32/S BUFX2
XFILL_51_DFFSR_239 INVX1_39/gnd DFFSR_54/S FILL
XFILL_14_3 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_27_DFFSR_138 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_16_XOR2X1_6 BUFX2_99/A DFFSR_7/S FILL
XFILL_9_OAI21X1_57 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_41_DFFSR_242 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_3_INVX1_185 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_26_DFFPOSX1_26 AND2X2_38/B DFFSR_23/S FILL
XFILL_47_DFFSR_93 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_17_DFFSR_141 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_3_CLKBUF1_6 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_1_NAND3X1_174 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_8_OAI21X1_60 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_31_DFFSR_245 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_21_DFFSR_248 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_8_AND2X2_2 BUFX2_99/A DFFSR_7/S FILL
XFILL_7_OAI21X1_63 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_6_NAND2X1_81 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_3_DFFSR_90 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_3_INVX1_37 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_31_DFFSR_43 BUFX2_98/A DFFSR_6/S FILL
XFILL_31_0_1 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_20_DFFSR_83 INVX1_3/gnd DFFSR_79/S FILL
XFILL_2_NOR2X1_20 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_6_DFFPOSX1_48 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_6_OAI21X1_66 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_5_NAND2X1_84 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_11_DFFSR_251 BUFX2_7/gnd DFFSR_151/S FILL
XNAND2X1_81 AND2X2_35/Y INVX1_143/Y DFFSR_34/gnd INVX1_157/A DFFSR_34/S NAND2X1
XFILL_4_NAND2X1_87 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_5_OAI21X1_69 INVX1_3/gnd DFFSR_23/S FILL
XOAI21X1_66 INVX1_160/A AND2X2_39/Y NAND2X1_85/Y XOR2X1_4/gnd OAI21X1_66/Y DFFSR_91/S
+ OAI21X1
XFILL_29_2_2 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_2_NAND3X1_108 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_3_DFFSR_138 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_3_NAND2X1_90 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_4_OAI21X1_72 INVX1_3/gnd DFFSR_23/S FILL
XFILL_2_BUFX2_28 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_44_DFFSR_169 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_2_NAND2X1_93 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_3_OAI21X1_75 INVX1_39/gnd DFFSR_54/S FILL
XFILL_1_DFFSR_3 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_7_DFFSR_245 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_4_NAND2X1_144 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_34_DFFSR_172 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_2_OAI21X1_78 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_1_NAND2X1_96 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_48_DFFSR_276 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_24_DFFSR_175 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_1_OAI21X1_81 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_0_NAND2X1_99 INVX1_39/gnd DFFSR_54/S FILL
XFILL_9_3_2 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_50_DFFSR_10 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_39_DFFSR_50 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_38_DFFSR_279 BUFX2_99/A DFFSR_7/S FILL
XFILL_0_INVX1_84 INVX1_39/gnd DFFSR_34/S FILL
XFILL_28_DFFSR_90 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_14_DFFSR_178 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_0_OAI21X1_84 BUFX2_98/A DFFSR_6/S FILL
XFILL_12_DFFSR_40 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_0_NAND3X1_204 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_1_OAI21X1_5 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_0_DFFSR_175 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_27_DFFSR_102 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_25_DFFSR_7 BUFX2_79/A DFFSR_7/S FILL
XFILL_9_OAI21X1_21 AND2X2_38/B DFFSR_59/S FILL
XFILL_41_DFFSR_206 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_3_INVX1_149 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_47_DFFSR_57 BUFX2_79/A DFFSR_6/S FILL
XFILL_36_DFFSR_97 INVX1_1/gnd DFFSR_97/S FILL
XFILL_6_AND2X2_16 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_17_DFFSR_105 INVX1_1/gnd DFFSR_53/S FILL
XFILL_8_OAI21X1_24 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_31_DFFSR_209 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_1_NAND3X1_138 INVX1_67/gnd DFFSR_201/S FILL
XFILL_21_DFFSR_212 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_7_OAI21X1_27 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_6_NAND2X1_45 INVX1_39/gnd DFFSR_34/S FILL
XFILL_20_DFFSR_47 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_3_DFFSR_54 INVX1_39/gnd DFFSR_54/S FILL
XFILL_6_DFFPOSX1_12 AND2X2_38/B DFFSR_23/S FILL
XFILL_3_NAND2X1_174 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_5_NAND2X1_48 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_6_OAI21X1_30 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_11_DFFSR_215 DFFSR_34/gnd DFFSR_1/S FILL
XNAND2X1_45 DFFSR_245/D NOR2X1_34/Y INVX1_39/gnd OAI21X1_13/C DFFSR_34/S NAND2X1
XFILL_4_NAND2X1_51 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_5_OAI21X1_33 INVX1_3/gnd DFFSR_79/S FILL
XOAI21X1_30 INVX1_138/A INVX1_139/A OAI21X1_30/C DFFSR_1/gnd AOI21X1_12/C DFFSR_81/S
+ OAI21X1
XFILL_3_DFFSR_102 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_3_NAND2X1_54 AND2X2_38/B DFFSR_59/S FILL
XFILL_4_OAI21X1_36 BUFX2_8/gnd DFFSR_51/S FILL
XDFFPOSX1_48 AND2X2_37/B CLKBUF1_45/Y NOR2X1_82/Y XOR2X1_4/gnd DFFSR_97/S DFFPOSX1
XFILL_44_DFFSR_133 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_46_DFFSR_3 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_15_DFFPOSX1_31 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_2_NAND2X1_57 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_3_OAI21X1_39 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_7_DFFSR_209 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_4_NAND2X1_108 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_34_DFFSR_136 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_2_OAI21X1_42 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_1_NAND2X1_60 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_48_DFFSR_240 INVX1_39/gnd DFFSR_34/S FILL
XFILL_24_DFFSR_139 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_0_NAND2X1_63 AND2X2_38/B DFFSR_59/S FILL
XFILL_1_OAI21X1_45 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_38_DFFSR_243 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_10_AOI22X1_11 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_0_INVX1_48 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_0_INVX1_186 BUFX2_79/A DFFSR_6/S FILL
XFILL_39_DFFSR_14 INVX1_1/gnd DFFSR_53/S FILL
XFILL_17_DFFSR_94 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_28_DFFSR_54 INVX1_39/gnd DFFSR_54/S FILL
XFILL_14_DFFSR_142 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_0_CLKBUF1_7 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_19_8 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_0_OAI21X1_48 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_28_DFFSR_246 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_36_3 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_18_DFFSR_249 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_25_DFFPOSX1_20 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_9_AOI22X1_14 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_0_NAND3X1_168 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_8_AOI22X1_17 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_1_INVX1_5 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_9_NAND3X1_223 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_7_AOI22X1_20 INVX1_39/gnd DFFSR_34/S FILL
XFILL_51_DFFSR_167 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_0_DFFSR_139 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_5_DFFPOSX1_42 INVX1_39/gnd DFFSR_34/S FILL
XDFFSR_249 BUFX2_90/A CLKBUF1_2/Y BUFX2_67/Y DFFSR_276/S INVX1_68/A BUFX2_72/gnd DFFSR_276/S
+ DFFSR
XFILL_6_AOI22X1_23 INVX1_39/gnd DFFSR_34/S FILL
XFILL_3_INVX1_113 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_41_DFFSR_170 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_36_DFFSR_61 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_47_DFFSR_21 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_5_AOI22X1_26 INVX1_1/gnd DFFSR_97/S FILL
XFILL_4_DFFSR_246 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_1_NAND3X1_102 INVX1_3/gnd DFFSR_23/S FILL
XFILL_31_DFFSR_173 XOR2X1_1/gnd DFFSR_208/S FILL
XAOI22X1_23 AOI22X1_23/A AOI22X1_23/B AOI21X1_21/A AOI21X1_21/B INVX1_39/gnd OAI21X1_53/A
+ DFFSR_34/S AOI22X1
XFILL_45_DFFSR_277 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_4_AOI22X1_29 INVX1_1/gnd DFFSR_53/S FILL
XFILL_21_DFFSR_176 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_35_DFFSR_280 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_3_DFFSR_18 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_20_DFFSR_11 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_3_NAND2X1_138 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_5_NAND2X1_12 INVX1_3/gnd DFFSR_79/S FILL
XFILL_11_DFFSR_179 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_4_NAND2X1_15 BUFX2_99/A DFFSR_92/S FILL
XFILL_7_XOR2X1_15 BUFX2_99/A DFFSR_7/S FILL
XFILL_6_NOR2X1_55 INVX1_39/gnd DFFSR_54/S FILL
XFILL_3_NAND2X1_18 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_8_OAI21X1_3 BUFX2_99/A DFFSR_92/S FILL
XDFFPOSX1_12 NOR3X1_1/A CLKBUF1_48/Y NOR2X1_64/Y AND2X2_38/B DFFSR_23/S DFFPOSX1
XFILL_12_DFFSR_1 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_2_NAND2X1_21 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_44_DFFSR_68 BUFX2_98/A DFFSR_6/S FILL
XFILL_7_DFFSR_173 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_24_DFFPOSX1_50 INVX1_1/gnd DFFSR_53/S FILL
XFILL_34_DFFSR_100 INVX1_1/gnd DFFSR_97/S FILL
XFILL_1_NAND2X1_24 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_48_DFFSR_204 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_24_DFFSR_103 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_8_NAND3X1_80 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_0_NAND2X1_27 AND2X2_38/B DFFSR_23/S FILL
XFILL_0_INVX1_12 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_0_DFFSR_65 BUFX2_79/A DFFSR_7/S FILL
XFILL_30_3_0 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_0_INVX1_150 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_38_DFFSR_207 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_17_DFFSR_58 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_3_AND2X2_17 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_28_DFFSR_18 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_14_DFFSR_106 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_7_NAND3X1_83 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_4_BUFX2_93 AND2X2_38/B DFFSR_59/S FILL
XFILL_28_DFFSR_210 BUFX2_98/A DFFSR_6/S FILL
XFILL_0_OAI21X1_12 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_6_NAND3X1_86 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_18_DFFSR_213 INVX1_3/gnd DFFSR_23/S FILL
XFILL_28_5_1 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_5_NAND3X1_89 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_0_NAND3X1_132 AND2X2_38/B DFFSR_23/S FILL
XNAND3X1_86 DFFSR_195/Q BUFX2_27/Y NOR2X1_31/Y DFFSR_62/gnd NAND3X1_86/Y DFFSR_62/S
+ NAND3X1
XFILL_4_NAND3X1_92 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_51_DFFSR_131 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_0_DFFSR_103 DFFSR_8/gnd DFFSR_60/S FILL
XDFFSR_213 INVX1_92/A CLKBUF1_12/Y BUFX2_70/Y DFFSR_23/S INVX1_93/A INVX1_3/gnd DFFSR_23/S
+ DFFSR
XFILL_3_NAND3X1_95 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_2_NAND2X1_168 BUFX2_79/A DFFSR_6/S FILL
XFILL_8_6_1 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_41_DFFSR_134 INVX1_1/gnd DFFSR_53/S FILL
XFILL_2_NAND3X1_98 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_8_DFFSR_72 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_36_DFFSR_25 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_25_DFFSR_65 BUFX2_79/A DFFSR_7/S FILL
XFILL_4_DFFSR_210 BUFX2_98/A DFFSR_6/S FILL
XFILL_31_DFFSR_137 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_45_DFFSR_241 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_7_CLKBUF1_5 BUFX2_99/A DFFSR_92/S FILL
XFILL_21_DFFSR_140 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_14_DFFPOSX1_25 BUFX2_79/A DFFSR_6/S FILL
XFILL_35_DFFSR_244 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_11_DFFSR_143 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_3_NAND2X1_102 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_25_DFFSR_247 BUFX2_99/A DFFSR_7/S FILL
XFILL_6_NOR2X1_19 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_15_DFFSR_250 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_11_OAI22X1_20 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_10_OAI22X1_23 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_44_DFFSR_32 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_7_DFFSR_137 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_33_DFFSR_72 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_24_DFFPOSX1_14 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_48_DFFSR_168 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_8_NAND3X1_44 BUFX2_99/A DFFSR_7/S FILL
XFILL_9_OAI22X1_26 INVX1_39/gnd DFFSR_54/S FILL
XFILL_0_INVX1_114 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_0_DFFSR_29 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_38_DFFSR_171 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_8_NAND3X1_217 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_17_DFFSR_22 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_7_NAND3X1_47 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_38_0_1 BUFX2_79/A DFFSR_7/S FILL
XFILL_1_DFFSR_247 BUFX2_99/A DFFSR_7/S FILL
XFILL_8_OAI22X1_29 INVX1_3/gnd DFFSR_79/S FILL
XFILL_4_BUFX2_57 AND2X2_38/B DFFSR_23/S FILL
XFILL_4_DFFPOSX1_36 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_28_DFFSR_174 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_42_DFFSR_278 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_6_NAND3X1_50 BUFX2_98/A DFFSR_6/S FILL
XFILL_7_OAI22X1_32 INVX1_39/gnd DFFSR_54/S FILL
XFILL_18_DFFSR_177 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_8_NOR3X1_3 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_5_NAND3X1_53 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_6_OAI22X1_35 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_36_2_2 BUFX2_99/A DFFSR_92/S FILL
XNAND3X1_50 DFFSR_7/Q NOR2X1_4/Y BUFX2_18/Y BUFX2_98/A AND2X2_12/B DFFSR_6/S NAND3X1
XFILL_4_NAND3X1_56 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_5_OAI22X1_38 AND2X2_38/B DFFSR_23/S FILL
XFILL_9_NAND3X1_151 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_41_DFFSR_79 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_3_NOR2X1_56 AND2X2_38/B DFFSR_59/S FILL
XOAI22X1_35 INVX1_85/Y OAI22X1_41/B INVX1_86/Y OAI22X1_41/D DFFSR_34/gnd NOR2X1_44/A
+ DFFSR_1/S OAI22X1
XFILL_3_NAND3X1_59 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_5_OAI21X1_4 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_4_OAI22X1_41 INVX1_39/gnd DFFSR_54/S FILL
XDFFSR_177 INVX1_60/A CLKBUF1_20/Y BUFX2_69/Y DFFSR_54/S INVX1_61/A DFFSR_46/gnd DFFSR_54/S
+ DFFSR
XFILL_2_NAND2X1_132 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_2_NAND3X1_62 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_3_OAI22X1_44 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_25_DFFSR_29 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_8_DFFSR_36 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_14_DFFSR_69 BUFX2_98/A DFFSR_32/S FILL
XFILL_4_DFFSR_174 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_31_DFFSR_101 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_2_OAI22X1_47 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_1_NAND3X1_65 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_45_DFFSR_205 INVX1_3/gnd DFFSR_79/S FILL
XFILL_0_NAND3X1_68 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_21_DFFSR_104 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_1_OAI22X1_50 INVX1_3/gnd DFFSR_23/S FILL
XFILL_0_OAI21X1_114 AND2X2_38/B DFFSR_59/S FILL
XFILL_35_DFFSR_208 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_0_AND2X2_18 AND2X2_38/B DFFSR_59/S FILL
XFILL_23_DFFPOSX1_44 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_11_DFFSR_107 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_25_DFFSR_211 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_1_XOR2X1_6 BUFX2_99/A DFFSR_7/S FILL
XFILL_49_DFFSR_86 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_15_DFFSR_214 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_7_NAND3X1_247 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_18_CLKBUF1_9 OR2X2_4/gnd DFFSR_3/S FILL
XINVX1_70 INVX1_70/A NOR3X1_6/gnd INVX1_70/Y DFFSR_79/S INVX1
XFILL_5_DFFSR_83 INVX1_3/gnd DFFSR_79/S FILL
XFILL_7_DFFSR_101 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_33_DFFSR_36 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_22_DFFSR_76 BUFX2_79/A DFFSR_7/S FILL
XFILL_48_DFFSR_132 INVX1_3/gnd DFFSR_79/S FILL
XINVX1_188 DFFSR_8/D BUFX2_77/gnd INVX1_188/Y DFFSR_98/S INVX1
XFILL_8_NAND3X1_181 INVX1_39/gnd DFFSR_54/S FILL
XFILL_38_DFFSR_135 DFFSR_62/gnd DFFSR_208/S FILL
XCLKBUF1_9 BUFX2_1/Y OR2X2_4/gnd DFFSR_7/CLK DFFSR_3/S CLKBUF1
XFILL_7_NAND3X1_11 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_1_DFFSR_211 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_4_BUFX2_21 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_28_DFFSR_138 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_1_NAND2X1_162 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_42_DFFSR_242 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_4_INVX1_185 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_6_NAND3X1_14 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_18_DFFSR_141 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_4_CLKBUF1_6 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_32_DFFSR_245 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_24_DFFSR_4 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_5_NAND3X1_17 BUFX2_99/A DFFSR_7/S FILL
XFILL_22_DFFSR_248 DFFSR_28/gnd DFFSR_8/S FILL
XNAND3X1_14 DFFSR_66/Q BUFX2_15/Y NOR2X1_2/Y DFFSR_4/gnd NAND3X1_14/Y DFFSR_4/S NAND3X1
XFILL_9_NAND3X1_115 BUFX2_79/A DFFSR_7/S FILL
XFILL_4_NAND3X1_20 BUFX2_99/A DFFSR_7/S FILL
XFILL_41_DFFSR_43 BUFX2_98/A DFFSR_6/S FILL
XFILL_30_DFFSR_83 INVX1_3/gnd DFFSR_79/S FILL
XFILL_2_INVX1_77 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_3_NOR2X1_20 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_13_DFFPOSX1_19 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_12_DFFSR_251 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_3_NAND3X1_23 OR2X2_6/gnd DFFSR_53/S FILL
XDFFSR_141 DFFSR_141/Q CLKBUF1_39/Y BUFX2_70/Y DFFSR_91/S INVX1_90/A XOR2X1_4/gnd
+ DFFSR_91/S DFFSR
XFILL_2_NAND3X1_26 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_14_DFFSR_33 BUFX2_98/A DFFSR_32/S FILL
XFILL_4_DFFSR_138 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_1_NAND3X1_29 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_2_OAI22X1_11 BUFX2_99/A DFFSR_92/S FILL
XFILL_1_BUFX2_68 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_45_DFFSR_169 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_0_NAND3X1_32 BUFX2_79/A DFFSR_7/S FILL
XFILL_1_OAI22X1_14 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_8_DFFSR_245 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_35_DFFSR_172 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_49_DFFSR_276 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_0_OAI22X1_17 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_25_DFFSR_175 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_49_DFFSR_50 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_39_DFFSR_279 BUFX2_99/A DFFSR_7/S FILL
XFILL_38_DFFSR_90 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_15_DFFSR_178 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_7_NAND3X1_211 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_3_DFFPOSX1_30 BUFX2_77/gnd DFFSR_98/S FILL
XDFFSR_87 INVX1_47/A CLKBUF1_38/Y DFFSR_15/R DFFSR_5/S DFFSR_79/Q BUFX2_77/gnd DFFSR_5/S
+ DFFSR
XFILL_5_DFFSR_47 BUFX2_77/gnd DFFSR_98/S FILL
XINVX1_34 DFFSR_77/Q OR2X2_4/gnd INVX1_34/Y DFFSR_3/S INVX1
XFILL_10_0_2 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_22_DFFSR_40 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_11_DFFSR_80 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_0_NOR2X1_57 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_2_OAI21X1_5 DFFSR_8/gnd DFFSR_8/S FILL
XINVX1_152 INVX1_152/A DFFSR_1/gnd INVX1_152/Y DFFSR_81/S INVX1
XFILL_8_NAND3X1_145 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_0_INVX1_2 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_1_4 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_1_DFFSR_175 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_12_DFFPOSX1_49 BUFX2_99/A DFFSR_92/S FILL
XFILL_28_DFFSR_102 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_42_DFFSR_206 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_1_NAND2X1_126 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_4_INVX1_149 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_46_DFFSR_97 INVX1_1/gnd DFFSR_97/S FILL
XFILL_7_AND2X2_16 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_18_DFFSR_105 INVX1_1/gnd DFFSR_53/S FILL
XFILL_32_DFFSR_209 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_22_DFFSR_212 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_7_AND2X2_6 BUFX2_99/A DFFSR_7/S FILL
XFILL_2_INVX1_41 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_30_DFFSR_47 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_2_DFFSR_94 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_19_DFFSR_87 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_12_DFFSR_215 DFFSR_34/gnd DFFSR_1/S FILL
XDFFSR_105 DFFSR_105/Q DFFSR_9/CLK BUFX2_49/Y DFFSR_53/S DFFSR_97/Q INVX1_1/gnd DFFSR_53/S
+ DFFSR
XFILL_22_DFFPOSX1_38 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_4_DFFSR_102 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_37_3_0 BUFX2_99/A DFFSR_7/S FILL
XFILL_6_NAND3X1_241 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_1_BUFX2_32 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_45_DFFSR_133 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_8_DFFSR_209 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_35_DFFSR_136 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_35_5_1 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_49_DFFSR_240 INVX1_39/gnd DFFSR_34/S FILL
XFILL_25_DFFSR_139 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_39_DFFSR_243 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_1_INVX1_186 BUFX2_79/A DFFSR_6/S FILL
XFILL_49_DFFSR_14 INVX1_1/gnd DFFSR_53/S FILL
XFILL_27_DFFSR_94 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_38_DFFSR_54 INVX1_39/gnd DFFSR_54/S FILL
XFILL_15_DFFSR_142 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_1_CLKBUF1_7 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_7_NAND3X1_175 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_29_DFFSR_246 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_0_NAND2X1_156 AND2X2_38/B DFFSR_59/S FILL
XFILL_19_DFFSR_249 BUFX2_72/gnd DFFSR_276/S FILL
XDFFSR_51 DFFSR_11/D CLKBUF1_8/Y DFFSR_1/R DFFSR_51/S DFFSR_51/D BUFX2_8/gnd DFFSR_51/S
+ DFFSR
XFILL_5_DFFSR_11 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_11_DFFSR_44 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_0_NOR2X1_21 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_8_NAND3X1_109 XOR2X1_1/gnd DFFSR_151/S FILL
XINVX1_116 DFFSR_160/Q DFFSR_5/gnd INVX1_116/Y DFFSR_5/S INVX1
XFILL_1_DFFSR_139 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_12_DFFPOSX1_13 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_4_INVX1_113 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_42_DFFSR_170 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_46_DFFSR_61 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_5_DFFSR_246 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_32_DFFSR_173 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_46_DFFSR_277 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_22_DFFSR_176 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_2_DFFSR_58 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_36_DFFSR_280 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_30_DFFSR_11 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_19_DFFSR_51 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_6_BUFX2_86 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_12_DFFSR_179 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_8_XOR2X1_15 BUFX2_99/A DFFSR_7/S FILL
XFILL_20_CLKBUF1_41 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_6_NAND3X1_205 INVX1_1/gnd DFFSR_53/S FILL
XFILL_45_0_1 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_36_DFFSR_7 BUFX2_79/A DFFSR_7/S FILL
XFILL_2_DFFPOSX1_24 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_19_CLKBUF1_44 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_8_DFFSR_173 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_35_DFFSR_100 INVX1_1/gnd DFFSR_97/S FILL
XAND2X2_20 AND2X2_20/A AND2X2_20/B OR2X2_6/gnd AND2X2_20/Y DFFSR_53/S AND2X2
XFILL_49_DFFSR_204 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_18_CLKBUF1_47 BUFX2_98/A DFFSR_32/S FILL
XFILL_25_DFFSR_103 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_43_2_2 OR2X2_4/gnd DFFSR_3/S FILL
XNAND3X1_241 INVX1_172/A AOI21X1_39/B AOI21X1_39/A DFFSR_8/gnd NAND3X1_243/B DFFSR_8/S
+ NAND3X1
XFILL_1_INVX1_150 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_39_DFFSR_207 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_27_DFFSR_58 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_16_DFFSR_98 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_4_AND2X2_17 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_38_DFFSR_18 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_15_DFFSR_106 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_7_NAND3X1_139 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_29_DFFSR_210 BUFX2_98/A DFFSR_6/S FILL
XFILL_11_DFFPOSX1_43 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_0_NAND2X1_120 DFFSR_46/gnd DFFSR_54/S FILL
XDFFSR_15 DFFSR_71/D CLKBUF1_37/Y DFFSR_15/R DFFSR_4/S DFFSR_15/D OR2X2_3/gnd DFFSR_4/S
+ DFFSR
XFILL_19_DFFSR_213 INVX1_3/gnd DFFSR_23/S FILL
XFILL_1_DFFSR_103 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_21_DFFPOSX1_32 INVX1_67/gnd DFFSR_201/S FILL
XFILL_42_DFFSR_134 INVX1_1/gnd DFFSR_53/S FILL
XFILL_11_1_0 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_46_DFFSR_25 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_35_DFFSR_65 BUFX2_79/A DFFSR_7/S FILL
XFILL_5_DFFSR_210 BUFX2_98/A DFFSR_6/S FILL
XFILL_32_DFFSR_137 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_46_DFFSR_241 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_5_NAND3X1_235 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_8_CLKBUF1_5 BUFX2_99/A DFFSR_92/S FILL
XFILL_22_DFFSR_140 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_2_DFFSR_22 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_36_DFFSR_244 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_19_DFFSR_15 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_12_DFFSR_143 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_6_BUFX2_50 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_26_DFFSR_247 BUFX2_99/A DFFSR_7/S FILL
XFILL_16_DFFSR_250 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_1_NOR2X1_3 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_6_NAND3X1_169 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_8_DFFSR_137 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_43_DFFSR_72 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_49_DFFSR_168 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_18_CLKBUF1_11 BUFX2_8/gnd DFFSR_51/S FILL
XNAND3X1_205 NAND3X1_203/A OAI21X1_67/Y AOI21X1_30/Y INVX1_1/gnd AOI22X1_29/C DFFSR_53/S
+ NAND3X1
XFILL_1_INVX1_114 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_39_DFFSR_171 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_17_CLKBUF1_14 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_27_DFFSR_22 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_16_DFFSR_62 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_2_DFFSR_247 BUFX2_99/A DFFSR_7/S FILL
XFILL_7_NAND3X1_103 AND2X2_38/B DFFSR_23/S FILL
XFILL_3_BUFX2_97 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_29_DFFSR_174 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_16_CLKBUF1_17 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_43_DFFSR_278 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_15_CLKBUF1_20 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_19_DFFSR_177 DFFSR_46/gnd DFFSR_54/S FILL
XNOR2X1_59 BUFX2_38/Y AOI21X1_1/A DFFSR_34/gnd NOR2X1_59/Y DFFSR_1/S NOR2X1
XFILL_14_CLKBUF1_23 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_13_CLKBUF1_26 INVX1_1/gnd DFFSR_53/S FILL
XFILL_4_NOR2X1_56 AND2X2_38/B DFFSR_59/S FILL
XFILL_23_DFFSR_1 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_6_OAI21X1_4 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_12_CLKBUF1_29 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_35_DFFSR_29 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_7_DFFSR_76 BUFX2_79/A DFFSR_7/S FILL
XFILL_24_DFFSR_69 BUFX2_98/A DFFSR_32/S FILL
XFILL_11_CLKBUF1_32 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_5_DFFSR_174 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_32_DFFSR_101 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_10_CLKBUF1_35 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_5_NAND3X1_199 INVX1_1/gnd DFFSR_97/S FILL
XFILL_46_DFFSR_205 INVX1_3/gnd DFFSR_79/S FILL
XFILL_22_DFFSR_104 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_1_DFFPOSX1_18 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_36_DFFSR_208 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_1_AND2X2_18 AND2X2_38/B DFFSR_59/S FILL
XFILL_17_0_2 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_6_BUFX2_14 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_12_DFFSR_107 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_26_DFFSR_211 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_9_CLKBUF1_38 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_16_DFFSR_214 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_8_CLKBUF1_41 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_6_NAND3X1_133 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_7_CLKBUF1_44 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_10_DFFPOSX1_37 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_19_CLKBUF1_9 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_8_DFFSR_101 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_43_DFFSR_36 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_32_DFFSR_76 BUFX2_79/A DFFSR_7/S FILL
XFILL_4_INVX1_70 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_6_CLKBUF1_47 BUFX2_98/A DFFSR_32/S FILL
XFILL_49_DFFSR_132 INVX1_3/gnd DFFSR_79/S FILL
XNAND3X1_169 INVX1_156/A OAI21X1_43/Y NAND2X1_80/Y XOR2X1_1/gnd NAND3X1_169/Y DFFSR_208/S
+ NAND3X1
XFILL_39_DFFSR_135 DFFSR_62/gnd DFFSR_208/S FILL
XCLKBUF1_47 clk BUFX2_98/A CLKBUF1_47/Y DFFSR_32/S CLKBUF1
XFILL_16_DFFSR_26 BUFX2_79/A DFFSR_6/S FILL
XFILL_2_DFFSR_211 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_3_BUFX2_61 AND2X2_38/B DFFSR_59/S FILL
XFILL_29_DFFSR_138 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_43_DFFSR_242 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_19_DFFSR_141 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_20_DFFPOSX1_26 AND2X2_38/B DFFSR_23/S FILL
XFILL_5_CLKBUF1_6 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_33_DFFSR_245 DFFSR_34/gnd DFFSR_34/S FILL
XNOR2X1_23 NOR2X1_23/A NOR2X1_23/B OR2X2_4/gnd NOR2X1_23/Y DFFSR_3/S NOR2X1
XFILL_44_3_0 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_23_DFFSR_248 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_4_NAND3X1_229 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_4_NOR2X1_20 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_40_DFFSR_83 INVX1_3/gnd DFFSR_79/S FILL
XFILL_13_DFFSR_251 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_0_DFFPOSX1_48 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_42_5_1 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_7_DFFSR_40 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_24_DFFSR_33 BUFX2_98/A DFFSR_32/S FILL
XFILL_13_DFFSR_73 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_5_DFFSR_138 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_5_NAND3X1_163 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_46_DFFSR_169 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_9_DFFSR_245 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_36_DFFSR_172 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_50_DFFSR_276 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_26_DFFSR_175 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_40_DFFSR_279 BUFX2_99/A DFFSR_7/S FILL
XFILL_48_DFFSR_90 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_16_DFFSR_178 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_32_DFFSR_40 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_21_DFFSR_80 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_4_DFFSR_87 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_4_INVX1_34 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_1_NOR2X1_57 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_6_CLKBUF1_11 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_3_OAI21X1_5 DFFSR_8/gnd DFFSR_8/S FILL
XNAND3X1_133 INVX1_127/Y INVX1_128/Y NOR2X1_61/Y BUFX2_8/gnd NAND3X1_134/B DFFSR_51/S
+ NAND3X1
XFILL_5_CLKBUF1_14 DFFSR_34/gnd DFFSR_34/S FILL
XCLKBUF1_11 BUFX2_4/Y BUFX2_8/gnd CLKBUF1_11/Y DFFSR_51/S CLKBUF1
XFILL_5_1 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_4_CLKBUF1_17 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_2_DFFSR_175 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_3_BUFX2_25 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_29_DFFSR_102 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_43_DFFSR_206 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_3_CLKBUF1_20 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_8_AND2X2_16 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_19_DFFSR_105 INVX1_1/gnd DFFSR_53/S FILL
XFILL_6_OAI21X1_115 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_33_DFFSR_209 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_14_DFFSR_8 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_2_CLKBUF1_23 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_13_NOR3X1_4 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_23_DFFSR_212 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_1_CLKBUF1_26 INVX1_1/gnd DFFSR_53/S FILL
XFILL_4_NAND3X1_193 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_1_INVX1_81 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_29_DFFSR_87 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_52_0_1 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_40_DFFSR_47 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_0_CLKBUF1_29 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_0_DFFPOSX1_12 AND2X2_38/B DFFSR_23/S FILL
XFILL_13_DFFSR_215 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_13_DFFSR_37 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_50_2_2 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_5_DFFSR_102 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_0_BUFX2_72 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_46_DFFSR_133 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_5_NAND3X1_127 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_9_DFFSR_209 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_36_DFFSR_136 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_50_DFFSR_240 INVX1_39/gnd DFFSR_34/S FILL
XFILL_35_DFFSR_4 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_26_DFFSR_139 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_40_DFFSR_243 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_37_DFFSR_94 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_2_INVX1_186 BUFX2_79/A DFFSR_6/S FILL
XFILL_48_DFFSR_54 INVX1_39/gnd DFFSR_54/S FILL
XFILL_16_DFFSR_142 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_2_CLKBUF1_7 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_30_DFFSR_246 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_20_DFFSR_249 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_21_DFFSR_44 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_4_DFFSR_51 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_1_NOR2X1_21 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_10_DFFSR_84 BUFX2_99/A DFFSR_7/S FILL
XFILL_18_1_0 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_19_DFFPOSX1_20 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_10_DFFSR_252 AND2X2_38/B DFFSR_23/S FILL
XFILL_3_NAND3X1_223 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_16_3_1 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_2_DFFSR_139 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_27_DFFPOSX1_8 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_43_DFFSR_170 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_6_DFFSR_246 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_33_DFFSR_173 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_14_5_2 INVX1_39/gnd DFFSR_54/S FILL
XFILL_47_DFFSR_277 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_23_DFFSR_176 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_4_NAND3X1_157 INVX1_3/gnd DFFSR_23/S FILL
XFILL_1_INVX1_45 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_37_DFFSR_280 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_40_DFFSR_11 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_1_DFFSR_98 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_18_DFFSR_91 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_29_DFFSR_51 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_13_DFFSR_179 OR2X2_1/gnd DFFSR_51/S FILL
XOAI21X1_115 XOR2X1_13/Y AOI21X1_67/A INVX1_212/Y NOR3X1_6/gnd AOI21X1_67/C DFFSR_91/S
+ OAI21X1
XFILL_9_DFFPOSX1_31 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_9_XOR2X1_15 BUFX2_99/A DFFSR_7/S FILL
XFILL_0_BUFX2_36 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_0_OAI21X1_6 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_9_DFFSR_173 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_36_DFFSR_100 INVX1_1/gnd DFFSR_97/S FILL
XFILL_18_DFFPOSX1_50 INVX1_1/gnd DFFSR_53/S FILL
XFILL_50_DFFSR_204 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_26_DFFSR_103 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_40_DFFSR_207 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_37_DFFSR_58 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_48_DFFSR_18 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_2_INVX1_150 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_26_DFFSR_98 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_5_AND2X2_17 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_16_DFFSR_106 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_30_DFFSR_210 BUFX2_98/A DFFSR_6/S FILL
XFILL_20_DFFSR_213 INVX1_3/gnd DFFSR_23/S FILL
XFILL_4_DFFSR_15 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_10_DFFSR_48 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_5_OAI21X1_109 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_10_DFFSR_216 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_3_NAND3X1_187 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_2_DFFSR_7 BUFX2_79/A DFFSR_7/S FILL
XFILL_2_DFFSR_103 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_24_0_2 AND2X2_38/B DFFSR_59/S FILL
XFILL_43_DFFSR_134 INVX1_1/gnd DFFSR_53/S FILL
XFILL_45_DFFSR_65 BUFX2_79/A DFFSR_7/S FILL
XFILL_6_DFFSR_210 BUFX2_98/A DFFSR_6/S FILL
XFILL_33_DFFSR_137 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_47_DFFSR_241 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_9_CLKBUF1_5 BUFX2_99/A DFFSR_92/S FILL
XFILL_23_DFFSR_140 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_4_NAND3X1_121 INVX1_1/gnd DFFSR_97/S FILL
XFILL_37_DFFSR_244 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_29_DFFSR_15 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_18_DFFSR_55 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_1_DFFSR_62 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_5_BUFX2_90 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_13_DFFSR_143 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_4_1_2 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_27_DFFSR_247 BUFX2_99/A DFFSR_7/S FILL
XFILL_6_NAND2X1_157 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_17_DFFSR_250 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_49_2 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_9_DFFSR_137 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_18_DFFPOSX1_14 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_50_DFFSR_168 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_40_DFFSR_171 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_51_3_0 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_2_INVX1_114 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_37_DFFSR_22 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_9_DFFSR_69 BUFX2_98/A DFFSR_32/S FILL
XFILL_26_DFFSR_62 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_2_NAND3X1_217 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_3_DFFSR_247 BUFX2_99/A DFFSR_7/S FILL
XFILL_30_DFFSR_174 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_44_DFFSR_278 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_17_DFFPOSX1_2 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_20_DFFSR_177 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_49_5_1 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_10_DFFSR_12 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_16_DFFPOSX1_5 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_10_DFFSR_180 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_15_DFFPOSX1_8 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_5_NOR2X1_56 AND2X2_38/B DFFSR_59/S FILL
XFILL_3_NAND3X1_151 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_47_DFFSR_7 BUFX2_79/A DFFSR_7/S FILL
XFILL_7_OAI21X1_4 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_8_DFFPOSX1_25 BUFX2_79/A DFFSR_6/S FILL
XFILL_45_DFFSR_29 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_34_DFFSR_69 BUFX2_98/A DFFSR_32/S FILL
XFILL_6_DFFSR_174 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_33_DFFSR_101 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_47_DFFSR_205 INVX1_3/gnd DFFSR_79/S FILL
XFILL_23_DFFSR_104 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_1_DFFSR_26 BUFX2_79/A DFFSR_6/S FILL
XFILL_37_DFFSR_208 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_18_DFFSR_19 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_2_AND2X2_18 AND2X2_38/B DFFSR_59/S FILL
XFILL_5_BUFX2_54 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_13_DFFSR_107 OR2X2_6/gnd DFFSR_92/S FILL
XBUFX2_94 BUFX2_94/A BUFX2_8/gnd BUFX2_94/Y DFFSR_51/S BUFX2
XFILL_17_DFFPOSX1_44 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_27_DFFSR_211 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_6_NAND2X1_121 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_2_INVX1_9 BUFX2_99/A DFFSR_7/S FILL
XFILL_17_DFFSR_214 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_15_6_0 INVX1_39/gnd DFFSR_34/S FILL
XFILL_0_NOR2X1_7 BUFX2_98/A DFFSR_32/S FILL
XFILL_1_NAND3X1_247 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_20_CLKBUF1_9 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_9_DFFSR_101 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_42_DFFSR_76 BUFX2_79/A DFFSR_7/S FILL
XNAND2X1_157 DFFSR_91/S NAND2X1_157/B NOR3X1_6/gnd AOI21X1_54/B DFFSR_91/S NAND2X1
XFILL_4_OAI21X1_103 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_50_DFFSR_132 INVX1_3/gnd DFFSR_79/S FILL
XFILL_8_AOI21X1_49 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_27_DFFPOSX1_33 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_40_DFFSR_135 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_9_DFFSR_33 BUFX2_98/A DFFSR_32/S FILL
XFILL_26_DFFSR_26 BUFX2_79/A DFFSR_6/S FILL
XFILL_7_AOI21X1_52 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_15_DFFSR_66 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_2_NAND3X1_181 INVX1_39/gnd DFFSR_54/S FILL
XFILL_3_DFFSR_211 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_30_DFFSR_138 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_44_DFFSR_242 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_6_AOI21X1_55 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_20_DFFSR_141 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_6_CLKBUF1_6 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_5_AOI21X1_58 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_34_DFFSR_245 DFFSR_34/gnd DFFSR_34/S FILL
XAOI21X1_55 AOI21X1_55/A AOI21X1_55/B NOR3X1_6/A XOR2X1_4/gnd AOI21X1_55/Y DFFSR_97/S
+ AOI21X1
XFILL_10_DFFSR_144 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_2_XOR2X1_3 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_4_AOI21X1_61 AND2X2_38/B DFFSR_59/S FILL
XFILL_24_DFFSR_248 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_5_NOR2X1_20 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_3_NAND3X1_115 BUFX2_79/A DFFSR_7/S FILL
XFILL_50_DFFSR_83 INVX1_3/gnd DFFSR_79/S FILL
XFILL_13_DFFSR_5 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_3_AOI21X1_64 AND2X2_38/B DFFSR_59/S FILL
XFILL_14_DFFSR_251 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_2_AOI21X1_67 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_54_7 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_5_NAND2X1_151 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_6_DFFSR_80 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_34_DFFSR_33 BUFX2_98/A DFFSR_32/S FILL
XFILL_23_DFFSR_73 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_1_AOI21X1_70 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_6_DFFSR_138 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_47_DFFSR_169 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_37_DFFSR_172 DFFSR_46/gnd DFFSR_62/S FILL
XBUFX2_58 BUFX2_58/A BUFX2_8/gnd BUFX2_58/Y DFFSR_81/S BUFX2
XFILL_0_DFFSR_248 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_5_BUFX2_18 BUFX2_98/A DFFSR_32/S FILL
XFILL_25_1_0 AND2X2_38/B DFFSR_23/S FILL
XFILL_27_DFFSR_175 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_9_OAI21X1_94 INVX1_67/gnd DFFSR_175/S FILL
XFILL_41_DFFSR_279 BUFX2_99/A DFFSR_7/S FILL
XFILL_17_DFFSR_178 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_8_OAI21X1_97 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_1_NAND3X1_211 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_34_DFFSR_1 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_23_3_1 OR2X2_1/gnd DFFSR_59/S FILL
XOAI21X1_8 INVX1_58/Y OAI21X1_4/B OAI21X1_8/C BUFX2_99/A OAI21X1_8/Y DFFSR_7/S OAI21X1
XFILL_42_DFFSR_40 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_3_INVX1_74 BUFX2_99/A DFFSR_92/S FILL
XFILL_31_DFFSR_80 DFFSR_4/gnd DFFSR_4/S FILL
XNAND2X1_121 DFFSR_3/S din[5] OR2X2_4/gnd OAI21X1_90/C DFFSR_32/S NAND2X1
XFILL_2_NOR2X1_57 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_5_2_0 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_4_OAI21X1_5 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_8_AOI21X1_13 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_21_5_2 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_7_AOI21X1_16 INVX1_67/gnd DFFSR_175/S FILL
XFILL_15_DFFSR_30 BUFX2_98/A DFFSR_32/S FILL
XFILL_2_NAND3X1_145 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_3_DFFSR_175 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_3_4_1 INVX1_67/gnd DFFSR_175/S FILL
XFILL_2_BUFX2_65 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_30_DFFSR_102 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_5_DFFPOSX1_2 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_6_AOI21X1_19 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_44_DFFSR_206 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_4_DFFPOSX1_5 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_20_DFFSR_105 INVX1_1/gnd DFFSR_53/S FILL
XFILL_7_DFFPOSX1_19 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_34_DFFSR_209 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_4_NAND2X1_181 BUFX2_99/A DFFSR_92/S FILL
XFILL_5_AOI21X1_22 DFFSR_62/gnd DFFSR_62/S FILL
XAOI21X1_19 NAND2X1_79/B OAI21X1_42/Y INVX1_154/A DFFSR_62/gnd AOI21X1_19/Y DFFSR_208/S
+ AOI21X1
XFILL_1_6_2 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_10_DFFSR_108 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_3_DFFPOSX1_8 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_4_AOI21X1_25 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_24_DFFSR_212 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_39_DFFSR_87 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_50_DFFSR_47 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_3_AOI21X1_28 AND2X2_38/B DFFSR_23/S FILL
XFILL_14_DFFSR_215 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_16_DFFPOSX1_38 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_2_AOI21X1_31 INVX1_39/gnd DFFSR_34/S FILL
XFILL_5_NAND2X1_115 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_23_DFFSR_37 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_6_DFFSR_44 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_12_DFFSR_77 BUFX2_98/A DFFSR_32/S FILL
XFILL_6_DFFSR_102 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_1_AOI21X1_34 INVX1_39/gnd DFFSR_34/S FILL
XFILL_0_NAND3X1_241 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_47_DFFSR_133 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_0_AOI21X1_37 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_37_DFFSR_136 NOR3X1_6/gnd DFFSR_79/S FILL
XBUFX2_22 AND2X2_4/Y OR2X2_6/gnd BUFX2_22/Y DFFSR_53/S BUFX2
XFILL_0_DFFSR_212 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_27_DFFSR_139 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_14_4 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_41_DFFSR_243 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_26_DFFPOSX1_27 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_9_OAI21X1_58 INVX1_39/gnd DFFSR_54/S FILL
XFILL_47_DFFSR_94 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_3_INVX1_186 BUFX2_79/A DFFSR_6/S FILL
XFILL_17_DFFSR_142 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_3_CLKBUF1_7 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_8_OAI21X1_61 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_1_NAND3X1_175 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_31_DFFSR_246 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_7_OAI21X1_64 INVX1_1/gnd DFFSR_53/S FILL
XFILL_6_NAND2X1_82 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_21_DFFSR_249 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_8_AND2X2_3 INVX1_1/gnd DFFSR_53/S FILL
XFILL_31_0_2 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_3_DFFSR_91 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_3_INVX1_38 AND2X2_38/B DFFSR_23/S FILL
XFILL_31_DFFSR_44 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_20_DFFSR_84 BUFX2_99/A DFFSR_7/S FILL
XFILL_6_DFFPOSX1_49 BUFX2_99/A DFFSR_92/S FILL
XFILL_2_NOR2X1_21 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_6_OAI21X1_67 INVX1_1/gnd DFFSR_97/S FILL
XFILL_5_NAND2X1_85 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_11_DFFSR_252 AND2X2_38/B DFFSR_23/S FILL
XNAND2X1_82 INVX1_133/A DFFSR_1/gnd DFFSR_1/gnd INVX1_158/A DFFSR_81/S NAND2X1
XFILL_5_OAI21X1_70 INVX1_3/gnd DFFSR_23/S FILL
XFILL_4_NAND2X1_88 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_2_NAND3X1_109 XOR2X1_1/gnd DFFSR_151/S FILL
XOAI21X1_67 INVX1_168/A NOR2X1_71/Y INVX1_167/Y INVX1_1/gnd OAI21X1_67/Y DFFSR_97/S
+ OAI21X1
XFILL_3_DFFSR_139 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_3_NAND2X1_91 INVX1_39/gnd DFFSR_54/S FILL
XFILL_4_OAI21X1_73 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_2_BUFX2_29 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_44_DFFSR_170 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_2_NAND2X1_94 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_3_OAI21X1_76 INVX1_1/gnd DFFSR_53/S FILL
XFILL_1_DFFSR_4 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_7_DFFSR_246 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_4_NAND2X1_145 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_34_DFFSR_173 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_48_DFFSR_277 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_2_OAI21X1_79 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_1_NAND2X1_97 INVX1_1/gnd DFFSR_97/S FILL
XFILL_24_DFFSR_176 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_1_OAI21X1_82 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_38_DFFSR_280 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_28_DFFSR_91 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_39_DFFSR_51 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_50_DFFSR_11 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_0_INVX1_85 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_14_DFFSR_179 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_0_OAI21X1_85 INVX1_39/gnd DFFSR_54/S FILL
XFILL_12_DFFSR_41 BUFX2_98/A DFFSR_6/S FILL
XFILL_1_OAI21X1_6 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_0_NAND3X1_205 INVX1_1/gnd DFFSR_53/S FILL
XFILL_37_DFFSR_100 INVX1_1/gnd DFFSR_97/S FILL
XFILL_0_DFFSR_176 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_27_DFFSR_103 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_25_DFFSR_8 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_41_DFFSR_207 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_47_DFFSR_58 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_3_INVX1_150 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_36_DFFSR_98 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_6_AND2X2_17 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_17_DFFSR_106 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_8_OAI21X1_25 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_31_DFFSR_210 BUFX2_98/A DFFSR_6/S FILL
XFILL_1_NAND3X1_139 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_7_OAI21X1_28 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_6_NAND2X1_46 INVX1_39/gnd DFFSR_34/S FILL
XFILL_21_DFFSR_213 INVX1_3/gnd DFFSR_23/S FILL
XFILL_3_DFFSR_55 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_20_DFFSR_48 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_6_DFFPOSX1_13 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_5_NAND2X1_49 INVX1_3/gnd DFFSR_79/S FILL
XFILL_11_DFFSR_216 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_3_NAND2X1_175 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_6_OAI21X1_31 AND2X2_38/B DFFSR_23/S FILL
XNAND2X1_46 DFFSR_165/Q AND2X2_18/Y INVX1_39/gnd NAND2X1_46/Y DFFSR_34/S NAND2X1
XFILL_5_OAI21X1_34 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_4_NAND2X1_52 OR2X2_6/gnd DFFSR_53/S FILL
XOAI21X1_31 INVX1_135/Y INVX1_145/Y OAI21X1_31/C AND2X2_38/B AOI22X1_19/C DFFSR_23/S
+ OAI21X1
XFILL_3_DFFSR_103 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_4_OAI21X1_37 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_3_NAND2X1_55 INVX1_39/gnd DFFSR_34/S FILL
XDFFPOSX1_49 AOI22X1_25/B CLKBUF1_46/Y AOI21X1_70/Y BUFX2_99/A DFFSR_92/S DFFPOSX1
XFILL_44_DFFSR_134 INVX1_1/gnd DFFSR_53/S FILL
XFILL_15_DFFPOSX1_32 INVX1_67/gnd DFFSR_201/S FILL
XFILL_2_NAND2X1_58 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_3_OAI21X1_40 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_46_DFFSR_4 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_7_DFFSR_210 BUFX2_98/A DFFSR_6/S FILL
XFILL_34_DFFSR_137 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_4_NAND2X1_109 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_48_DFFSR_241 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_1_NAND2X1_61 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_2_OAI21X1_43 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_22_6_0 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_24_DFFSR_140 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_1_OAI21X1_46 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_0_NAND2X1_64 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_39_DFFSR_15 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_28_DFFSR_55 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_0_INVX1_49 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_0_INVX1_187 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_38_DFFSR_244 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_10_AOI22X1_12 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_17_DFFSR_95 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_14_DFFSR_143 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_0_CLKBUF1_8 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_19_9 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_0_OAI21X1_49 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_28_DFFSR_247 BUFX2_99/A DFFSR_7/S FILL
XFILL_36_4 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_25_DFFPOSX1_21 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_18_DFFSR_250 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_9_AOI22X1_15 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_8_AOI22X1_18 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_1_INVX1_6 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_0_NAND3X1_169 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_7_AOI22X1_21 AND2X2_38/B DFFSR_59/S FILL
XFILL_5_DFFPOSX1_43 OR2X2_2/gnd DFFSR_216/S FILL
XDFFSR_250 BUFX2_91/A DFFSR_85/CLK BUFX2_65/Y DFFSR_8/S INVX1_75/A DFFSR_8/gnd DFFSR_8/S
+ DFFSR
XFILL_0_DFFSR_140 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_6_AOI22X1_24 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_41_DFFSR_171 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_3_INVX1_114 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_47_DFFSR_22 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_36_DFFSR_62 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_4_DFFSR_247 BUFX2_99/A DFFSR_7/S FILL
XFILL_5_AOI22X1_27 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_1_NAND3X1_103 AND2X2_38/B DFFSR_23/S FILL
XFILL_31_DFFSR_174 BUFX2_8/gnd DFFSR_51/S FILL
XAOI22X1_24 AOI22X1_24/A AOI22X1_24/B AOI21X1_22/A AOI21X1_22/B DFFSR_46/gnd OAI21X1_53/B
+ DFFSR_62/S AOI22X1
XFILL_45_DFFSR_278 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_6_NAND2X1_10 BUFX2_79/A DFFSR_7/S FILL
XFILL_21_DFFSR_177 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_3_DFFSR_19 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_20_DFFSR_12 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_5_NAND2X1_13 BUFX2_99/A DFFSR_92/S FILL
XFILL_3_NAND2X1_139 INVX1_1/gnd DFFSR_97/S FILL
XFILL_11_DFFSR_180 DFFSR_34/gnd DFFSR_34/S FILL
XNAND2X1_10 AND2X2_3/Y NOR2X1_1/Y BUFX2_79/A OAI21X1_4/B DFFSR_7/S NAND2X1
XFILL_4_NAND2X1_16 BUFX2_79/A DFFSR_7/S FILL
XFILL_6_NOR2X1_56 AND2X2_38/B DFFSR_59/S FILL
XFILL_8_OAI21X1_4 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_3_NAND2X1_19 DFFSR_8/gnd DFFSR_8/S FILL
XDFFPOSX1_13 INVX1_3/A CLKBUF1_43/Y AOI21X1_6/Y BUFX2_8/gnd DFFSR_81/S DFFPOSX1
XFILL_12_DFFSR_2 BUFX2_79/A DFFSR_7/S FILL
XFILL_2_NAND2X1_22 BUFX2_99/A DFFSR_7/S FILL
XFILL_32_1_0 INVX1_1/gnd DFFSR_97/S FILL
XFILL_44_DFFSR_69 BUFX2_98/A DFFSR_32/S FILL
XFILL_7_DFFSR_174 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_34_DFFSR_101 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_9_NAND3X1_78 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_1_NAND2X1_25 BUFX2_99/A DFFSR_7/S FILL
XFILL_48_DFFSR_205 INVX1_3/gnd DFFSR_79/S FILL
XFILL_24_DFFSR_104 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_8_NAND3X1_81 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_1_OAI21X1_10 BUFX2_79/A DFFSR_7/S FILL
XFILL_30_3_1 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_0_NAND2X1_28 AND2X2_38/B DFFSR_59/S FILL
XFILL_38_DFFSR_208 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_28_DFFSR_19 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_0_INVX1_13 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_0_DFFSR_66 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_0_INVX1_151 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_17_DFFSR_59 AND2X2_38/B DFFSR_59/S FILL
XFILL_3_AND2X2_18 AND2X2_38/B DFFSR_59/S FILL
XFILL_14_DFFSR_107 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_7_NAND3X1_84 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_4_BUFX2_94 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_0_OAI21X1_13 INVX1_39/gnd DFFSR_54/S FILL
XFILL_28_DFFSR_211 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_6_NAND3X1_87 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_18_DFFSR_214 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_28_5_2 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_5_NAND3X1_90 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_0_NAND3X1_133 BUFX2_8/gnd DFFSR_51/S FILL
XNAND3X1_87 NAND3X1_87/A NAND3X1_86/Y AOI22X1_11/Y DFFSR_46/gnd NOR2X1_43/B DFFSR_62/S
+ NAND3X1
XFILL_21_CLKBUF1_9 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_9_NAND3X1_188 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_4_NAND3X1_93 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_3_NAND3X1_96 DFFSR_34/gnd DFFSR_1/S FILL
XDFFSR_214 INVX1_99/A CLKBUF1_25/Y BUFX2_60/Y DFFSR_276/S DFFSR_214/D BUFX2_72/gnd
+ DFFSR_276/S DFFSR
XFILL_0_DFFSR_104 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_2_NAND2X1_169 INVX1_1/gnd DFFSR_53/S FILL
XFILL_8_6_2 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_41_DFFSR_135 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_8_DFFSR_73 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_2_NAND3X1_99 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_25_DFFSR_66 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_36_DFFSR_26 BUFX2_79/A DFFSR_6/S FILL
XFILL_4_DFFSR_211 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_31_DFFSR_138 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_45_DFFSR_242 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_21_DFFSR_141 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_7_CLKBUF1_6 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_14_DFFPOSX1_26 AND2X2_38/B DFFSR_23/S FILL
XFILL_35_DFFSR_245 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_7_BUFX2_11 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_3_NAND2X1_103 AND2X2_38/B DFFSR_23/S FILL
XFILL_11_DFFSR_144 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_25_DFFSR_248 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_6_NOR2X1_20 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_15_DFFSR_251 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_11_OAI22X1_21 BUFX2_98/A DFFSR_32/S FILL
XFILL_10_OAI22X1_24 BUFX2_98/A DFFSR_32/S FILL
XFILL_44_DFFSR_33 BUFX2_98/A DFFSR_32/S FILL
XFILL_33_DFFSR_73 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_7_DFFSR_138 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_24_DFFPOSX1_15 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_9_NAND3X1_42 BUFX2_79/A DFFSR_6/S FILL
XFILL_48_DFFSR_169 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_9_OAI22X1_27 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_8_NAND3X1_45 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_38_DFFSR_172 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_0_DFFSR_30 BUFX2_98/A DFFSR_32/S FILL
XFILL_0_INVX1_115 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_17_DFFSR_23 AND2X2_38/B DFFSR_23/S FILL
XFILL_8_NAND3X1_218 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_7_NAND3X1_48 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_1_DFFSR_248 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_38_0_2 BUFX2_79/A DFFSR_7/S FILL
XFILL_8_OAI22X1_30 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_4_BUFX2_58 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_4_DFFPOSX1_37 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_28_DFFSR_175 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_42_DFFSR_279 BUFX2_99/A DFFSR_7/S FILL
XFILL_6_NAND3X1_51 BUFX2_99/A DFFSR_7/S FILL
XFILL_7_OAI22X1_33 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_18_DFFSR_178 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_8_NOR3X1_4 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_6_OAI22X1_36 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_5_NAND3X1_54 OR2X2_3/gnd DFFSR_60/S FILL
XNAND3X1_51 BUFX2_88/A AND2X2_3/Y BUFX2_22/Y BUFX2_99/A AND2X2_12/A DFFSR_7/S NAND3X1
XFILL_4_NAND3X1_57 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_5_OAI22X1_39 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_41_DFFSR_80 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_3_NOR2X1_57 XOR2X1_4/gnd DFFSR_91/S FILL
XOAI22X1_36 INVX1_87/Y OAI22X1_45/B INVX1_88/Y OAI22X1_45/D BUFX2_7/gnd NOR2X1_45/A
+ DFFSR_216/S OAI22X1
XFILL_5_OAI21X1_5 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_3_NAND3X1_60 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_4_OAI22X1_42 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_2_NAND2X1_133 BUFX2_72/gnd DFFSR_201/S FILL
XDFFSR_178 INVX1_69/A CLKBUF1_12/Y BUFX2_70/Y DFFSR_79/S INVX1_70/A NOR3X1_6/gnd DFFSR_79/S
+ DFFSR
XFILL_3_OAI22X1_45 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_2_NAND3X1_63 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_8_DFFSR_37 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_14_DFFSR_70 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_25_DFFSR_30 BUFX2_98/A DFFSR_32/S FILL
XFILL_4_DFFSR_175 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_31_DFFSR_102 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_1_NAND3X1_66 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_2_OAI22X1_48 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_45_DFFSR_206 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_0_NAND3X1_69 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_21_DFFSR_105 INVX1_1/gnd DFFSR_53/S FILL
XFILL_1_OAI22X1_51 INVX1_39/gnd DFFSR_54/S FILL
XFILL_35_DFFSR_209 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_0_OAI21X1_115 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_0_AND2X2_19 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_23_DFFPOSX1_45 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_11_DFFSR_108 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_25_DFFSR_212 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_1_XOR2X1_7 BUFX2_98/A DFFSR_6/S FILL
XFILL_0_DFFSR_1 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_49_DFFSR_87 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_7_NAND3X1_248 INVX1_3/gnd DFFSR_79/S FILL
XFILL_15_DFFSR_215 DFFSR_34/gnd DFFSR_1/S FILL
XINVX1_71 INVX1_71/A BUFX2_79/A INVX1_71/Y DFFSR_6/S INVX1
XFILL_33_DFFSR_37 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_5_DFFSR_84 BUFX2_99/A DFFSR_7/S FILL
XFILL_7_DFFSR_102 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_22_DFFSR_77 BUFX2_98/A DFFSR_32/S FILL
XFILL_48_DFFSR_133 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_38_DFFSR_136 NOR3X1_6/gnd DFFSR_79/S FILL
XINVX1_189 NOR3X1_6/A XOR2X1_4/gnd DFFSR_257/R DFFSR_91/S INVX1
XFILL_8_NAND3X1_182 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_1_DFFSR_212 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_7_NAND3X1_12 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_18_1 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_4_BUFX2_22 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_28_DFFSR_139 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_1_NAND2X1_163 INVX1_67/gnd DFFSR_201/S FILL
XFILL_42_DFFSR_243 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_6_NAND3X1_15 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_4_INVX1_186 BUFX2_79/A DFFSR_6/S FILL
XFILL_18_DFFSR_142 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_4_CLKBUF1_7 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_24_DFFSR_5 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_14_NOR3X1_1 INVX1_3/gnd DFFSR_79/S FILL
XFILL_32_DFFSR_246 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_5_NAND3X1_18 BUFX2_79/A DFFSR_7/S FILL
XNAND3X1_15 NAND3X1_13/Y NAND3X1_14/Y AOI22X1_2/Y DFFSR_4/gnd NOR2X1_11/B DFFSR_4/S
+ NAND3X1
XFILL_22_DFFSR_249 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_4_NAND3X1_21 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_41_DFFSR_44 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_30_DFFSR_84 BUFX2_99/A DFFSR_7/S FILL
XFILL_2_INVX1_78 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_3_NOR2X1_21 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_12_DFFSR_252 AND2X2_38/B DFFSR_23/S FILL
XFILL_13_DFFPOSX1_20 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_3_NAND3X1_24 INVX1_1/gnd DFFSR_97/S FILL
XDFFSR_142 DFFSR_198/D CLKBUF1_15/Y BUFX2_60/Y DFFSR_151/S INVX1_97/A XOR2X1_1/gnd
+ DFFSR_151/S DFFSR
XFILL_2_NAND3X1_27 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_29_6_0 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_14_DFFSR_34 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_4_DFFSR_139 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_1_BUFX2_69 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_2_OAI22X1_12 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_1_NAND3X1_30 BUFX2_79/A DFFSR_6/S FILL
XFILL_45_DFFSR_170 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_1_OAI22X1_15 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_0_NAND3X1_33 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_8_DFFSR_246 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_35_DFFSR_173 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_49_DFFSR_277 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_0_OAI22X1_18 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_45_DFFSR_1 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_25_DFFSR_176 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_39_DFFSR_280 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_38_DFFSR_91 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_49_DFFSR_51 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_15_DFFSR_179 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_7_NAND3X1_212 INVX1_39/gnd DFFSR_54/S FILL
XFILL_3_DFFPOSX1_31 XOR2X1_4/gnd DFFSR_97/S FILL
XINVX1_35 INVX1_35/A DFFSR_28/gnd INVX1_35/Y DFFSR_3/S INVX1
XDFFSR_88 INVX1_54/A DFFSR_85/CLK DFFSR_5/R DFFSR_98/S DFFSR_80/Q DFFSR_4/gnd DFFSR_98/S
+ DFFSR
XFILL_5_DFFSR_48 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_22_DFFSR_41 BUFX2_98/A DFFSR_6/S FILL
XFILL_11_DFFSR_81 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_0_NOR2X1_58 INVX1_3/gnd DFFSR_79/S FILL
XFILL_2_OAI21X1_6 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_38_DFFSR_100 INVX1_1/gnd DFFSR_97/S FILL
XINVX1_153 INVX1_153/A INVX1_67/gnd INVX1_153/Y DFFSR_175/S INVX1
XFILL_8_NAND3X1_146 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_1_5 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_1_DFFSR_176 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_0_INVX1_3 INVX1_3/gnd DFFSR_79/S FILL
XFILL_12_DFFPOSX1_50 INVX1_1/gnd DFFSR_53/S FILL
XFILL_28_DFFSR_103 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_1_NAND2X1_127 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_42_DFFSR_207 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_4_INVX1_150 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_46_DFFSR_98 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_7_AND2X2_17 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_18_DFFSR_106 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_32_DFFSR_210 BUFX2_98/A DFFSR_6/S FILL
XFILL_7_AND2X2_7 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_22_DFFSR_213 INVX1_3/gnd DFFSR_23/S FILL
XFILL_30_DFFSR_48 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_19_DFFSR_88 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_2_DFFSR_95 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_2_INVX1_42 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_39_1_0 BUFX2_79/A DFFSR_6/S FILL
XFILL_12_DFFSR_216 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_22_DFFPOSX1_39 BUFX2_7/gnd DFFSR_151/S FILL
XDFFSR_106 DFFSR_114/D CLKBUF1_27/Y BUFX2_49/Y DFFSR_91/S DFFSR_98/Q XOR2X1_4/gnd
+ DFFSR_91/S DFFSR
XFILL_4_DFFSR_103 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_37_3_1 BUFX2_99/A DFFSR_7/S FILL
XFILL_6_NAND3X1_242 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_1_BUFX2_33 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_45_DFFSR_134 INVX1_1/gnd DFFSR_53/S FILL
XFILL_8_DFFSR_210 BUFX2_98/A DFFSR_6/S FILL
XFILL_35_DFFSR_137 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_49_DFFSR_241 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_35_5_2 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_25_DFFSR_140 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_49_DFFSR_15 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_38_DFFSR_55 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_1_INVX1_187 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_39_DFFSR_244 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_27_DFFSR_95 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_15_DFFSR_143 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_7_NAND3X1_176 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_1_CLKBUF1_8 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_29_DFFSR_247 BUFX2_99/A DFFSR_7/S FILL
XFILL_19_DFFSR_250 DFFSR_8/gnd DFFSR_8/S FILL
XDFFSR_52 DFFSR_12/D CLKBUF1_4/Y DFFSR_8/R DFFSR_4/S INVX1_25/A OR2X2_3/gnd DFFSR_4/S
+ DFFSR
XFILL_0_NAND2X1_157 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_5_DFFSR_12 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_11_DFFSR_45 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_0_NOR2X1_22 OR2X2_4/gnd DFFSR_3/S FILL
XINVX1_117 INVX1_117/A BUFX2_7/gnd INVX1_117/Y DFFSR_151/S INVX1
XFILL_8_NAND3X1_110 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_1_DFFSR_140 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_12_DFFPOSX1_14 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_42_DFFSR_171 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_4_INVX1_114 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_46_DFFSR_62 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_5_DFFSR_247 BUFX2_99/A DFFSR_7/S FILL
XFILL_32_DFFSR_174 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_46_DFFSR_278 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_22_DFFSR_177 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_30_DFFSR_12 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_19_DFFSR_52 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_2_DFFSR_59 AND2X2_38/B DFFSR_59/S FILL
XFILL_6_BUFX2_87 INVX1_1/gnd DFFSR_53/S FILL
XFILL_12_DFFSR_180 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_9_OAI21X1_4 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_20_CLKBUF1_42 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_6_NAND3X1_206 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_45_0_2 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_36_DFFSR_8 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_2_DFFPOSX1_25 BUFX2_79/A DFFSR_6/S FILL
XFILL_19_CLKBUF1_45 BUFX2_79/A DFFSR_7/S FILL
XFILL_8_DFFSR_174 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_35_DFFSR_101 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_18_CLKBUF1_48 INVX1_3/gnd DFFSR_79/S FILL
XFILL_49_DFFSR_205 INVX1_3/gnd DFFSR_79/S FILL
XAND2X2_21 AND2X2_21/A AND2X2_21/B DFFSR_34/gnd AND2X2_21/Y DFFSR_34/S AND2X2
XNAND3X1_242 XOR2X1_8/B AOI21X1_38/B AOI21X1_38/A DFFSR_28/gnd NAND3X1_242/Y DFFSR_3/S
+ NAND3X1
XFILL_25_DFFSR_104 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_38_DFFSR_19 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_1_INVX1_151 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_39_DFFSR_208 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_16_DFFSR_99 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_27_DFFSR_59 AND2X2_38/B DFFSR_59/S FILL
XFILL_4_AND2X2_18 AND2X2_38/B DFFSR_59/S FILL
XFILL_15_DFFSR_107 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_7_NAND3X1_140 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_29_DFFSR_211 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_11_DFFPOSX1_44 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_19_DFFSR_214 BUFX2_72/gnd DFFSR_276/S FILL
XDFFSR_16 DFFSR_16/Q DFFSR_7/CLK DFFSR_9/R DFFSR_3/S DFFSR_16/D DFFSR_28/gnd DFFSR_3/S
+ DFFSR
XFILL_0_NAND2X1_121 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_1_DFFSR_104 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_21_DFFPOSX1_33 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_42_DFFSR_135 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_11_1_1 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_35_DFFSR_66 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_46_DFFSR_26 BUFX2_79/A DFFSR_6/S FILL
XFILL_5_DFFSR_211 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_32_DFFSR_138 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_46_DFFSR_242 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_5_NAND3X1_236 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_22_DFFSR_141 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_8_CLKBUF1_6 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_19_DFFSR_16 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_2_DFFSR_23 AND2X2_38/B DFFSR_23/S FILL
XFILL_36_DFFSR_245 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_6_BUFX2_51 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_12_DFFSR_144 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_26_DFFSR_248 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_16_DFFSR_251 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_1_NOR2X1_4 INVX1_1/gnd DFFSR_53/S FILL
XFILL_6_NAND3X1_170 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_43_DFFSR_73 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_8_DFFSR_138 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_18_CLKBUF1_12 AND2X2_38/B DFFSR_23/S FILL
XFILL_49_DFFSR_169 DFFSR_62/gnd DFFSR_62/S FILL
XNAND3X1_206 OAI21X1_69/Y INVX1_164/Y OAI21X1_70/Y BUFX2_8/gnd NAND3X1_214/B DFFSR_81/S
+ NAND3X1
XFILL_1_INVX1_115 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_17_CLKBUF1_15 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_39_DFFSR_172 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_16_DFFSR_63 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_27_DFFSR_23 AND2X2_38/B DFFSR_23/S FILL
XFILL_2_DFFSR_248 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_7_NAND3X1_104 AND2X2_38/B DFFSR_23/S FILL
XFILL_3_BUFX2_98 BUFX2_79/A DFFSR_7/S FILL
XFILL_29_DFFSR_175 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_16_CLKBUF1_18 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_43_DFFSR_279 BUFX2_99/A DFFSR_7/S FILL
XFILL_15_CLKBUF1_21 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_19_DFFSR_178 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_36_6_0 BUFX2_99/A DFFSR_92/S FILL
XNOR2X1_60 OR2X2_1/Y NOR2X1_60/B DFFSR_34/gnd NOR2X1_60/Y DFFSR_34/S NOR2X1
XFILL_14_CLKBUF1_24 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_23_DFFSR_2 BUFX2_79/A DFFSR_7/S FILL
XFILL_13_CLKBUF1_27 INVX1_1/gnd DFFSR_97/S FILL
XFILL_4_NOR2X1_57 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_6_OAI21X1_5 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_12_CLKBUF1_30 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_24_DFFSR_70 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_35_DFFSR_30 BUFX2_98/A DFFSR_32/S FILL
XFILL_7_DFFSR_77 BUFX2_98/A DFFSR_32/S FILL
XFILL_11_CLKBUF1_33 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_5_DFFSR_175 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_32_DFFSR_102 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_46_DFFSR_206 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_5_NAND3X1_200 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_10_CLKBUF1_36 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_22_DFFSR_105 INVX1_1/gnd DFFSR_53/S FILL
XFILL_36_DFFSR_209 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_1_DFFPOSX1_19 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_1_AND2X2_19 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_6_BUFX2_15 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_12_DFFSR_108 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_26_DFFSR_212 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_9_CLKBUF1_39 INVX1_1/gnd DFFSR_53/S FILL
XFILL_16_DFFSR_215 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_8_CLKBUF1_42 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_6_NAND3X1_134 INVX1_39/gnd DFFSR_54/S FILL
XFILL_7_CLKBUF1_45 BUFX2_79/A DFFSR_7/S FILL
XFILL_10_DFFPOSX1_38 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_43_DFFSR_37 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_4_INVX1_71 BUFX2_79/A DFFSR_6/S FILL
XFILL_8_DFFSR_102 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_32_DFFSR_77 BUFX2_98/A DFFSR_32/S FILL
XFILL_6_CLKBUF1_48 INVX1_3/gnd DFFSR_79/S FILL
XFILL_49_DFFSR_133 BUFX2_77/gnd DFFSR_5/S FILL
XNAND3X1_170 INVX1_131/Y NAND3X1_169/Y OAI21X1_44/Y XOR2X1_1/gnd OAI21X1_45/C DFFSR_208/S
+ NAND3X1
XFILL_39_DFFSR_136 NOR3X1_6/gnd DFFSR_79/S FILL
XCLKBUF1_48 clk INVX1_3/gnd CLKBUF1_48/Y DFFSR_79/S CLKBUF1
XFILL_16_DFFSR_27 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_2_DFFSR_212 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_3_BUFX2_62 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_46_1_0 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_29_DFFSR_139 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_43_DFFSR_243 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_19_DFFSR_142 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_5_CLKBUF1_7 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_20_DFFPOSX1_27 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_33_DFFSR_246 XOR2X1_1/gnd DFFSR_208/S FILL
XNOR2X1_24 NOR2X1_24/A NOR2X1_24/B DFFSR_4/gnd NOR2X1_24/Y DFFSR_4/S NOR2X1
XFILL_23_DFFSR_249 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_44_3_1 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_4_NAND3X1_230 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_40_DFFSR_84 BUFX2_99/A DFFSR_7/S FILL
XFILL_4_NOR2X1_21 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_0_DFFPOSX1_49 BUFX2_99/A DFFSR_92/S FILL
XFILL_13_DFFSR_252 AND2X2_38/B DFFSR_23/S FILL
XFILL_42_5_2 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_7_DFFSR_41 BUFX2_98/A DFFSR_6/S FILL
XFILL_24_DFFSR_34 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_13_DFFSR_74 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_5_DFFSR_139 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_46_DFFSR_170 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_5_NAND3X1_164 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_9_DFFSR_246 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_36_DFFSR_173 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_50_DFFSR_277 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_26_DFFSR_176 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_40_DFFSR_280 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_48_DFFSR_91 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_16_DFFSR_179 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_10_4_0 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_4_INVX1_35 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_4_DFFSR_88 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_32_DFFSR_41 BUFX2_98/A DFFSR_6/S FILL
XFILL_21_DFFSR_81 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_1_NOR2X1_58 INVX1_3/gnd DFFSR_79/S FILL
XFILL_6_CLKBUF1_12 AND2X2_38/B DFFSR_23/S FILL
XFILL_3_OAI21X1_6 OR2X2_4/gnd DFFSR_3/S FILL
XNAND3X1_134 INVX1_124/Y NAND3X1_134/B NAND2X1_55/Y INVX1_39/gnd DFFPOSX1_9/D DFFSR_54/S
+ NAND3X1
XFILL_5_CLKBUF1_15 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_39_DFFSR_100 INVX1_1/gnd DFFSR_97/S FILL
XCLKBUF1_12 BUFX2_5/Y AND2X2_38/B CLKBUF1_12/Y DFFSR_23/S CLKBUF1
XFILL_5_2 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_2_DFFSR_176 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_4_CLKBUF1_18 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_3_BUFX2_26 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_29_DFFSR_103 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_3_CLKBUF1_21 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_43_DFFSR_207 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_8_AND2X2_17 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_6_OAI21X1_116 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_19_DFFSR_106 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_2_CLKBUF1_24 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_33_DFFSR_210 BUFX2_98/A DFFSR_6/S FILL
XFILL_13_NOR3X1_5 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_14_DFFSR_9 BUFX2_79/A DFFSR_6/S FILL
XFILL_23_DFFSR_213 INVX1_3/gnd DFFSR_23/S FILL
XFILL_1_CLKBUF1_27 INVX1_1/gnd DFFSR_97/S FILL
XFILL_4_NAND3X1_194 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_1_INVX1_82 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_40_DFFSR_48 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_29_DFFSR_88 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_52_0_2 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_13_DFFSR_216 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_0_CLKBUF1_30 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_0_DFFPOSX1_13 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_5_DFFSR_103 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_13_DFFSR_38 BUFX2_98/A DFFSR_6/S FILL
XFILL_0_BUFX2_73 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_46_DFFSR_134 INVX1_1/gnd DFFSR_53/S FILL
XFILL_5_NAND3X1_128 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_9_DFFSR_210 BUFX2_98/A DFFSR_6/S FILL
XFILL_36_DFFSR_137 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_50_DFFSR_241 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_35_DFFSR_5 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_26_DFFSR_140 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_2_INVX1_187 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_40_DFFSR_244 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_48_DFFSR_55 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_37_DFFSR_95 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_16_DFFSR_143 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_2_CLKBUF1_8 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_30_DFFSR_247 BUFX2_99/A DFFSR_7/S FILL
XFILL_20_DFFSR_250 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_4_DFFSR_52 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_19_DFFPOSX1_21 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_10_DFFSR_85 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_21_DFFSR_45 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_1_NOR2X1_22 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_18_1_1 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_10_DFFSR_253 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_0_0_0 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_3_NAND3X1_224 INVX1_39/gnd DFFSR_54/S FILL
XFILL_16_3_2 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_2_DFFSR_140 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_27_DFFPOSX1_9 INVX1_67/gnd DFFSR_201/S FILL
XFILL_43_DFFSR_171 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_6_DFFSR_247 BUFX2_99/A DFFSR_7/S FILL
XFILL_33_DFFSR_174 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_47_DFFSR_278 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_4_NAND3X1_158 AND2X2_38/B DFFSR_59/S FILL
XFILL_23_DFFSR_177 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_40_DFFSR_12 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_29_DFFSR_52 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_1_INVX1_46 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_1_DFFSR_99 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_18_DFFSR_92 BUFX2_99/A DFFSR_92/S FILL
XFILL_13_DFFSR_180 DFFSR_34/gnd DFFSR_34/S FILL
XOAI21X1_116 NOR2X1_81/A NOR2X1_81/B OAI21X1_116/C XOR2X1_4/gnd OAI21X1_116/Y DFFSR_91/S
+ OAI21X1
XFILL_9_DFFPOSX1_32 INVX1_67/gnd DFFSR_201/S FILL
XFILL_0_BUFX2_37 INVX1_1/gnd DFFSR_97/S FILL
XFILL_0_OAI21X1_7 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_9_DFFSR_174 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_36_DFFSR_101 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_50_DFFSR_205 INVX1_3/gnd DFFSR_79/S FILL
XFILL_26_DFFSR_104 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_43_6_0 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_48_DFFSR_19 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_2_INVX1_151 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_40_DFFSR_208 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_26_DFFSR_99 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_37_DFFSR_59 AND2X2_38/B DFFSR_59/S FILL
XFILL_5_AND2X2_18 AND2X2_38/B DFFSR_59/S FILL
XFILL_16_DFFSR_107 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_30_DFFSR_211 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_20_DFFSR_214 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_4_DFFSR_16 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_10_DFFSR_49 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_5_OAI21X1_110 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_10_DFFSR_217 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_3_NAND3X1_188 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_2_DFFSR_104 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_2_DFFSR_8 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_43_DFFSR_135 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_45_DFFSR_66 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_6_DFFSR_211 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_33_DFFSR_138 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_47_DFFSR_242 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_4_NAND3X1_122 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_23_DFFSR_141 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_9_CLKBUF1_6 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_29_DFFSR_16 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_1_DFFSR_63 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_1_INVX1_10 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_37_DFFSR_245 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_18_DFFSR_56 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_13_DFFSR_144 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_5_BUFX2_91 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_27_DFFSR_248 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_6_NAND2X1_158 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_49_3 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_17_DFFSR_251 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_53_1_0 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_9_DFFSR_138 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_18_DFFPOSX1_15 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_50_DFFSR_169 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_2_INVX1_115 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_40_DFFSR_172 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_9_DFFSR_70 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_51_3_1 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_26_DFFSR_63 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_37_DFFSR_23 AND2X2_38/B DFFSR_23/S FILL
XFILL_2_NAND3X1_218 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_3_DFFSR_248 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_30_DFFSR_175 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_44_DFFSR_279 BUFX2_99/A DFFSR_7/S FILL
XFILL_17_DFFPOSX1_3 INVX1_39/gnd DFFSR_34/S FILL
XFILL_20_DFFSR_178 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_49_5_2 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_10_DFFSR_13 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_16_DFFPOSX1_6 AND2X2_38/B DFFSR_23/S FILL
XFILL_10_DFFSR_181 INVX1_3/gnd DFFSR_79/S FILL
XFILL_15_DFFPOSX1_9 INVX1_67/gnd DFFSR_201/S FILL
XFILL_5_NOR2X1_57 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_3_NAND3X1_152 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_47_DFFSR_8 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_7_OAI21X1_5 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_8_DFFPOSX1_26 AND2X2_38/B DFFSR_23/S FILL
XFILL_45_DFFSR_30 BUFX2_98/A DFFSR_32/S FILL
XFILL_6_DFFSR_175 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_34_DFFSR_70 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_33_DFFSR_102 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_47_DFFSR_206 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_23_DFFSR_105 INVX1_1/gnd DFFSR_53/S FILL
XFILL_37_DFFSR_209 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_1_DFFSR_27 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_2_AND2X2_19 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_18_DFFSR_20 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_17_4_0 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_13_DFFSR_108 OR2X2_6/gnd DFFSR_92/S FILL
XBUFX2_95 BUFX2_95/A BUFX2_8/gnd BUFX2_95/Y DFFSR_81/S BUFX2
XFILL_5_BUFX2_55 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_27_DFFSR_212 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_17_DFFPOSX1_45 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_10_OAI22X1_1 INVX1_1/gnd DFFSR_53/S FILL
XFILL_6_NAND2X1_122 INVX1_67/gnd DFFSR_175/S FILL
XFILL_17_DFFSR_215 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_9_NOR3X1_1 INVX1_3/gnd DFFSR_79/S FILL
XFILL_15_6_1 INVX1_39/gnd DFFSR_34/S FILL
XFILL_0_NOR2X1_8 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_1_NAND3X1_248 INVX1_3/gnd DFFSR_79/S FILL
XFILL_9_AOI21X1_47 INVX1_67/gnd DFFSR_175/S FILL
XFILL_9_DFFSR_102 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_42_DFFSR_77 BUFX2_98/A DFFSR_32/S FILL
XNAND2X1_158 NAND2X1_157/B INVX1_208/Y XOR2X1_4/gnd AOI21X1_55/A DFFSR_97/S NAND2X1
XFILL_50_DFFSR_133 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_4_OAI21X1_104 INVX1_67/gnd DFFSR_201/S FILL
XFILL_8_AOI21X1_50 INVX1_67/gnd DFFSR_175/S FILL
XFILL_27_DFFPOSX1_34 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_40_DFFSR_136 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_9_DFFSR_34 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_26_DFFSR_27 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_7_AOI21X1_53 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_15_DFFSR_67 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_2_NAND3X1_182 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_3_DFFSR_212 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_30_DFFSR_139 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_6_AOI21X1_56 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_44_DFFSR_243 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_20_DFFSR_142 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_6_CLKBUF1_7 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_5_AOI21X1_59 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_34_DFFSR_246 XOR2X1_1/gnd DFFSR_208/S FILL
XAOI21X1_56 AOI21X1_56/A AOI21X1_56/B NOR3X1_6/A NOR3X1_6/gnd AOI21X1_56/Y DFFSR_79/S
+ AOI21X1
XFILL_10_DFFSR_145 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_24_DFFSR_249 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_2_XOR2X1_4 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_4_AOI21X1_62 INVX1_3/gnd DFFSR_23/S FILL
XFILL_50_DFFSR_84 BUFX2_99/A DFFSR_7/S FILL
XFILL_5_NOR2X1_21 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_13_DFFSR_6 BUFX2_79/A DFFSR_6/S FILL
XFILL_3_NAND3X1_116 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_3_AOI21X1_65 INVX1_3/gnd DFFSR_23/S FILL
XFILL_14_DFFSR_252 AND2X2_38/B DFFSR_23/S FILL
XFILL_2_AOI21X1_68 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_54_8 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_5_NAND2X1_152 INVX1_1/gnd DFFSR_97/S FILL
XFILL_6_DFFSR_81 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_34_DFFSR_34 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_23_DFFSR_74 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_6_DFFSR_139 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_1_AOI21X1_71 BUFX2_99/A DFFSR_92/S FILL
XFILL_47_DFFSR_170 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_37_DFFSR_173 XOR2X1_1/gnd DFFSR_208/S FILL
XBUFX2_59 BUFX2_58/A AND2X2_38/B BUFX2_59/Y DFFSR_23/S BUFX2
XFILL_0_DFFSR_249 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_5_BUFX2_19 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_27_DFFSR_176 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_25_1_1 AND2X2_38/B DFFSR_23/S FILL
XFILL_9_OAI21X1_95 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_41_DFFSR_280 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_17_DFFSR_179 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_7_0_0 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_34_DFFSR_2 BUFX2_79/A DFFSR_7/S FILL
XFILL_8_OAI21X1_98 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_1_NAND3X1_212 INVX1_39/gnd DFFSR_54/S FILL
XFILL_23_3_2 OR2X2_1/gnd DFFSR_59/S FILL
XOAI21X1_9 INVX1_68/Y OAI21X1_9/B OAI21X1_9/C INVX1_67/gnd OAI21X1_9/Y DFFSR_201/S
+ OAI21X1
XFILL_42_DFFSR_41 BUFX2_98/A DFFSR_6/S FILL
XFILL_3_INVX1_75 BUFX2_98/A DFFSR_6/S FILL
XFILL_9_AOI21X1_11 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_31_DFFSR_81 DFFSR_1/gnd DFFSR_81/S FILL
XNAND2X1_122 DFFSR_276/S din[6] INVX1_67/gnd OAI21X1_91/C DFFSR_175/S NAND2X1
XFILL_2_NOR2X1_58 INVX1_3/gnd DFFSR_79/S FILL
XFILL_5_2_1 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_4_OAI21X1_6 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_8_AOI21X1_14 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_40_DFFSR_100 INVX1_1/gnd DFFSR_97/S FILL
XFILL_7_AOI21X1_17 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_15_DFFSR_31 BUFX2_79/A DFFSR_6/S FILL
XFILL_3_DFFSR_176 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_2_NAND3X1_146 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_3_4_2 INVX1_67/gnd DFFSR_175/S FILL
XFILL_30_DFFSR_103 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_2_BUFX2_66 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_6_AOI21X1_20 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_5_DFFPOSX1_3 INVX1_39/gnd DFFSR_34/S FILL
XFILL_44_DFFSR_207 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_20_DFFSR_106 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_7_DFFPOSX1_20 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_4_DFFPOSX1_6 AND2X2_38/B DFFSR_23/S FILL
XFILL_5_AOI21X1_23 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_34_DFFSR_210 BUFX2_98/A DFFSR_6/S FILL
XFILL_4_NAND2X1_182 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_10_DFFSR_109 DFFSR_4/gnd DFFSR_4/S FILL
XAOI21X1_20 INVX1_152/Y AOI21X1_20/B OAI21X1_41/B DFFSR_1/gnd OAI21X1_53/C DFFSR_1/S
+ AOI21X1
XFILL_3_DFFPOSX1_9 INVX1_67/gnd DFFSR_201/S FILL
XFILL_24_DFFSR_213 INVX1_3/gnd DFFSR_23/S FILL
XFILL_4_AOI21X1_26 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_50_DFFSR_48 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_39_DFFSR_88 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_3_AOI21X1_29 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_14_DFFSR_216 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_16_DFFPOSX1_39 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_2_AOI21X1_32 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_6_DFFSR_45 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_50_6_0 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_5_NAND2X1_116 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_6_DFFSR_103 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_12_DFFSR_78 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_23_DFFSR_38 BUFX2_98/A DFFSR_6/S FILL
XFILL_1_AOI21X1_35 INVX1_39/gnd DFFSR_54/S FILL
XFILL_0_NAND3X1_242 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_47_DFFSR_134 INVX1_1/gnd DFFSR_53/S FILL
XFILL_0_AOI21X1_38 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_37_DFFSR_137 BUFX2_7/gnd DFFSR_216/S FILL
XBUFX2_23 BUFX2_23/A XOR2X1_1/gnd BUFX2_23/Y DFFSR_151/S BUFX2
XFILL_0_DFFSR_213 INVX1_3/gnd DFFSR_23/S FILL
XFILL_14_5 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_27_DFFSR_140 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_26_DFFPOSX1_28 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_3_INVX1_187 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_41_DFFSR_244 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_47_DFFSR_95 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_17_DFFSR_143 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_3_CLKBUF1_8 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_31_DFFSR_247 BUFX2_99/A DFFSR_7/S FILL
XFILL_8_OAI21X1_62 INVX1_3/gnd DFFSR_79/S FILL
XFILL_1_NAND3X1_176 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_7_OAI21X1_65 INVX1_1/gnd DFFSR_53/S FILL
XFILL_8_AND2X2_4 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_6_NAND2X1_83 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_21_DFFSR_250 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_20_DFFSR_85 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_31_DFFSR_45 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_3_DFFSR_92 BUFX2_99/A DFFSR_92/S FILL
XFILL_3_INVX1_39 INVX1_39/gnd DFFSR_34/S FILL
XFILL_2_NOR2X1_22 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_6_DFFPOSX1_50 INVX1_1/gnd DFFSR_53/S FILL
XFILL_6_OAI21X1_68 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_5_NAND2X1_86 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_11_DFFSR_253 DFFSR_34/gnd DFFSR_1/S FILL
XNAND2X1_83 AND2X2_35/Y AND2X2_36/Y DFFSR_34/gnd NAND2X1_83/Y DFFSR_34/S NAND2X1
XFILL_4_NAND2X1_89 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_5_OAI21X1_71 INVX1_3/gnd DFFSR_79/S FILL
XOAI21X1_68 INVX1_134/Y NOR2X1_69/B XOR2X1_4/Y OR2X2_6/gnd AOI22X1_28/A DFFSR_92/S
+ OAI21X1
XFILL_2_NAND3X1_110 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_3_DFFSR_140 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_3_NAND2X1_92 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_2_BUFX2_30 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_4_OAI21X1_74 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_44_DFFSR_171 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_3_OAI21X1_77 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_2_NAND2X1_95 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_1_DFFSR_5 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_7_DFFSR_247 BUFX2_99/A DFFSR_7/S FILL
XFILL_4_NAND2X1_146 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_34_DFFSR_174 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_2_OAI21X1_80 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_1_NAND2X1_98 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_48_DFFSR_278 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_24_DFFSR_177 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_50_DFFSR_12 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_1_OAI21X1_83 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_39_DFFSR_52 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_28_DFFSR_92 BUFX2_99/A DFFSR_92/S FILL
XFILL_0_INVX1_86 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_14_DFFSR_180 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_0_OAI21X1_86 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_12_DFFSR_42 OR2X2_4/gnd DFFSR_32/S FILL
XBUFX2_1 BUFX2_3/A OR2X2_4/gnd BUFX2_1/Y DFFSR_32/S BUFX2
XFILL_0_NAND3X1_206 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_1_OAI21X1_7 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_37_DFFSR_101 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_51_DFFSR_205 INVX1_3/gnd DFFSR_79/S FILL
XFILL_0_DFFSR_177 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_27_DFFSR_104 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_25_DFFSR_9 BUFX2_79/A DFFSR_6/S FILL
XFILL_3_INVX1_151 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_41_DFFSR_208 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_36_DFFSR_99 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_47_DFFSR_59 AND2X2_38/B DFFSR_59/S FILL
XFILL_6_AND2X2_18 AND2X2_38/B DFFSR_59/S FILL
XFILL_17_DFFSR_107 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_8_OAI21X1_26 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_31_DFFSR_211 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_1_NAND3X1_140 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_21_DFFSR_214 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_7_OAI21X1_29 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_6_NAND2X1_47 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_3_DFFSR_56 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_20_DFFSR_49 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_6_DFFPOSX1_14 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_3_NAND2X1_176 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_6_OAI21X1_32 AND2X2_38/B DFFSR_59/S FILL
XFILL_5_NAND2X1_50 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_11_DFFSR_217 BUFX2_72/gnd DFFSR_201/S FILL
XNAND2X1_47 DFFSR_238/Q NOR2X1_34/Y DFFSR_62/gnd NAND2X1_47/Y DFFSR_208/S NAND2X1
XFILL_4_NAND2X1_53 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_5_OAI21X1_35 BUFX2_7/gnd DFFSR_216/S FILL
XOAI21X1_32 INVX1_135/Y INVX1_145/Y AND2X2_32/Y AND2X2_38/B OAI21X1_32/Y DFFSR_59/S
+ OAI21X1
XFILL_3_DFFSR_104 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_3_NAND2X1_56 AND2X2_38/B DFFSR_59/S FILL
XFILL_4_OAI21X1_38 OR2X2_1/gnd DFFSR_59/S FILL
XDFFPOSX1_50 DFFPOSX1_50/Q CLKBUF1_45/Y NOR2X1_83/Y INVX1_1/gnd DFFSR_53/S DFFPOSX1
XFILL_24_4_0 AND2X2_38/B DFFSR_59/S FILL
XFILL_44_DFFSR_135 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_46_DFFSR_5 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_15_DFFPOSX1_33 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_3_OAI21X1_41 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_2_NAND2X1_59 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_7_DFFSR_211 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_4_NAND2X1_110 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_34_DFFSR_138 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_1_NAND2X1_62 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_2_OAI21X1_44 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_48_DFFSR_242 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_22_6_1 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_24_DFFSR_141 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_0_NAND2X1_65 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_0_INVX1_50 BUFX2_98/A DFFSR_6/S FILL
XFILL_1_OAI21X1_47 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_38_DFFSR_245 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_39_DFFSR_16 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_28_DFFSR_56 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_17_DFFSR_96 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_0_INVX1_188 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_10_AOI22X1_13 AND2X2_38/B DFFSR_23/S FILL
XFILL_4_5_0 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_0_CLKBUF1_9 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_14_DFFSR_144 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_28_DFFSR_248 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_0_OAI21X1_50 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_36_5 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_18_DFFSR_251 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_9_AOI22X1_16 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_25_DFFPOSX1_22 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_0_NAND3X1_170 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_1_INVX1_7 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_8_AOI22X1_19 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_9_NAND3X1_225 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_7_AOI22X1_22 INVX1_3/gnd DFFSR_79/S FILL
XFILL_5_DFFPOSX1_44 OR2X2_2/gnd DFFSR_216/S FILL
XDFFSR_251 BUFX2_92/A CLKBUF1_20/Y BUFX2_62/Y DFFSR_151/S INVX1_82/A BUFX2_7/gnd DFFSR_151/S
+ DFFSR
XFILL_0_DFFSR_141 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_6_AOI22X1_25 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_3_INVX1_115 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_41_DFFSR_172 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_36_DFFSR_63 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_47_DFFSR_23 AND2X2_38/B DFFSR_23/S FILL
XFILL_4_DFFSR_248 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_5_AOI22X1_28 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_31_DFFSR_175 OR2X2_2/gnd DFFSR_175/S FILL
XAOI22X1_25 BUFX2_59/Y AOI22X1_25/B INVX1_135/A AND2X2_37/B XOR2X1_4/gnd INVX1_168/A
+ DFFSR_97/S AOI22X1
XFILL_1_NAND3X1_104 AND2X2_38/B DFFSR_23/S FILL
XFILL_45_DFFSR_279 BUFX2_99/A DFFSR_7/S FILL
XFILL_6_NAND2X1_11 BUFX2_98/A DFFSR_6/S FILL
XFILL_21_DFFSR_178 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_3_DFFSR_20 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_20_DFFSR_13 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_3_NAND2X1_140 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_5_NAND2X1_14 BUFX2_98/A DFFSR_32/S FILL
XFILL_11_DFFSR_181 INVX1_3/gnd DFFSR_79/S FILL
XNAND2X1_11 DFFSR_41/D AND2X2_5/Y BUFX2_98/A NAND3X1_4/A DFFSR_6/S NAND2X1
XFILL_4_NAND2X1_17 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_6_NOR2X1_57 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_8_OAI21X1_5 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_2_NOR2X1_1 BUFX2_99/A DFFSR_92/S FILL
XFILL_3_NAND2X1_20 DFFSR_8/gnd DFFSR_8/S FILL
XDFFPOSX1_14 NAND2X1_59/A CLKBUF1_47/Y XOR2X1_1/Y DFFSR_62/gnd DFFSR_62/S DFFPOSX1
XFILL_12_DFFSR_3 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_2_NAND2X1_23 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_32_1_1 INVX1_1/gnd DFFSR_97/S FILL
XFILL_7_DFFSR_175 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_44_DFFSR_70 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_34_DFFSR_102 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_9_NAND3X1_79 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_1_NAND2X1_26 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_48_DFFSR_206 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_24_DFFSR_105 INVX1_1/gnd DFFSR_53/S FILL
XFILL_0_NAND2X1_29 INVX1_3/gnd DFFSR_23/S FILL
XFILL_8_NAND3X1_82 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_38_DFFSR_209 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_0_INVX1_14 BUFX2_98/A DFFSR_6/S FILL
XFILL_30_3_2 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_0_INVX1_152 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_1_OAI21X1_11 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_3_AND2X2_19 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_17_DFFSR_60 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_28_DFFSR_20 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_0_DFFSR_67 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_14_DFFSR_108 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_4_BUFX2_95 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_7_NAND3X1_85 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_28_DFFSR_212 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_0_OAI21X1_14 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_6_NAND3X1_88 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_18_DFFSR_215 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_5_NAND3X1_91 AND2X2_38/B DFFSR_59/S FILL
XFILL_0_NAND3X1_134 INVX1_39/gnd DFFSR_54/S FILL
XNAND3X1_88 NOR2X1_41/Y NOR2X1_42/Y NOR2X1_43/Y DFFSR_1/gnd XOR2X1_10/B DFFSR_81/S
+ NAND3X1
XFILL_4_NAND3X1_94 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_0_DFFSR_105 INVX1_1/gnd DFFSR_53/S FILL
XFILL_3_NAND3X1_97 AND2X2_38/B DFFSR_59/S FILL
XFILL_2_NAND2X1_170 BUFX2_7/gnd DFFSR_216/S FILL
XDFFSR_215 INVX1_106/A CLKBUF1_29/Y BUFX2_66/Y DFFSR_1/S DFFSR_207/Q DFFSR_34/gnd
+ DFFSR_1/S DFFSR
XFILL_41_DFFSR_136 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_36_DFFSR_27 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_8_DFFSR_74 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_25_DFFSR_67 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_4_DFFSR_212 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_31_DFFSR_139 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_45_DFFSR_243 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_21_DFFSR_142 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_7_CLKBUF1_7 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_14_DFFPOSX1_27 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_35_DFFSR_246 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_3_NAND2X1_104 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_11_DFFSR_145 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_25_DFFSR_249 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_6_NOR2X1_21 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_15_DFFSR_252 AND2X2_38/B DFFSR_23/S FILL
XFILL_10_OAI22X1_25 INVX1_39/gnd DFFSR_54/S FILL
XFILL_33_DFFSR_74 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_44_DFFSR_34 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_7_DFFSR_139 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_24_DFFPOSX1_16 INVX1_67/gnd DFFSR_175/S FILL
XFILL_48_DFFSR_170 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_8_NAND3X1_46 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_9_OAI22X1_28 INVX1_3/gnd DFFSR_23/S FILL
XFILL_0_INVX1_116 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_0_DFFSR_31 BUFX2_79/A DFFSR_6/S FILL
XFILL_8_NAND3X1_219 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_38_DFFSR_173 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_17_DFFSR_24 BUFX2_98/A DFFSR_6/S FILL
XFILL_1_DFFSR_249 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_7_NAND3X1_49 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_4_BUFX2_59 AND2X2_38/B DFFSR_23/S FILL
XFILL_8_OAI22X1_31 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_28_DFFSR_176 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_4_DFFPOSX1_38 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_42_DFFSR_280 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_6_NAND3X1_52 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_7_OAI22X1_34 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_18_DFFSR_179 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_8_NOR3X1_5 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_5_NAND3X1_55 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_6_OAI22X1_37 INVX1_3/gnd DFFSR_23/S FILL
XNAND3X1_52 NAND3X1_52/A NAND3X1_49/Y AND2X2_12/Y DFFSR_8/gnd NOR2X1_26/A DFFSR_60/S
+ NAND3X1
XFILL_4_NAND3X1_58 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_41_DFFSR_81 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_5_OAI22X1_40 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_3_NOR2X1_58 INVX1_3/gnd DFFSR_79/S FILL
XOAI22X1_37 INVX1_90/Y OAI22X1_43/B INVX1_91/Y OAI22X1_43/D INVX1_3/gnd NOR2X1_47/B
+ DFFSR_23/S OAI22X1
XFILL_3_NAND3X1_61 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_5_OAI21X1_6 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_4_OAI22X1_43 DFFSR_62/gnd DFFSR_208/S FILL
XDFFSR_179 INVX1_76/A CLKBUF1_22/Y BUFX2_61/Y DFFSR_51/S INVX1_77/A OR2X2_1/gnd DFFSR_51/S
+ DFFSR
XFILL_2_NAND2X1_134 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_2_NAND3X1_64 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_41_DFFSR_100 INVX1_1/gnd DFFSR_97/S FILL
XFILL_3_OAI22X1_46 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_8_DFFSR_38 BUFX2_98/A DFFSR_6/S FILL
XFILL_25_DFFSR_31 BUFX2_79/A DFFSR_6/S FILL
XFILL_14_DFFSR_71 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_4_DFFSR_176 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_1_NAND3X1_67 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_31_DFFSR_103 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_2_OAI22X1_49 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_45_DFFSR_207 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_21_DFFSR_106 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_0_NAND3X1_70 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_1_OAI22X1_52 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_35_DFFSR_210 BUFX2_98/A DFFSR_6/S FILL
XFILL_0_OAI21X1_116 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_0_AND2X2_20 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_23_DFFPOSX1_46 INVX1_39/gnd DFFSR_34/S FILL
XFILL_11_DFFSR_109 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_1_XOR2X1_8 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_0_DFFSR_2 BUFX2_79/A DFFSR_7/S FILL
XFILL_25_DFFSR_213 INVX1_3/gnd DFFSR_23/S FILL
XFILL_49_DFFSR_88 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_15_DFFSR_216 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_7_NAND3X1_249 OR2X2_6/gnd DFFSR_92/S FILL
XINVX1_72 INVX1_72/A NOR3X1_6/gnd INVX1_72/Y DFFSR_79/S INVX1
XFILL_5_DFFSR_85 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_7_DFFSR_103 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_22_DFFSR_78 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_33_DFFSR_38 BUFX2_98/A DFFSR_6/S FILL
XFILL_48_DFFSR_134 INVX1_1/gnd DFFSR_53/S FILL
XFILL_8_NAND3X1_10 BUFX2_79/A DFFSR_6/S FILL
XFILL_38_DFFSR_137 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_8_NAND3X1_183 OR2X2_1/gnd DFFSR_59/S FILL
XINVX1_190 DFFSR_265/Q OR2X2_2/gnd INVX1_190/Y DFFSR_216/S INVX1
XFILL_18_2 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_4_BUFX2_23 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_7_NAND3X1_13 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_1_DFFSR_213 INVX1_3/gnd DFFSR_23/S FILL
XFILL_28_DFFSR_140 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_1_NAND2X1_164 INVX1_67/gnd DFFSR_175/S FILL
XFILL_42_DFFSR_244 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_6_NAND3X1_16 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_4_INVX1_187 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_4_CLKBUF1_8 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_18_DFFSR_143 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_32_DFFSR_247 BUFX2_99/A DFFSR_7/S FILL
XFILL_24_DFFSR_6 BUFX2_79/A DFFSR_6/S FILL
XFILL_5_NAND3X1_19 BUFX2_99/A DFFSR_92/S FILL
XFILL_14_NOR3X1_2 INVX1_1/gnd DFFSR_53/S FILL
XNAND3X1_16 NOR2X1_9/Y NOR2X1_10/Y NOR2X1_11/Y DFFSR_28/gnd XOR2X1_9/A DFFSR_8/S NAND3X1
XFILL_22_DFFSR_250 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_31_4_0 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_9_NAND3X1_117 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_41_DFFSR_45 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_4_NAND3X1_22 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_2_INVX1_79 INVX1_39/gnd DFFSR_54/S FILL
XFILL_3_NOR2X1_22 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_30_DFFSR_85 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_13_DFFPOSX1_21 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_12_DFFSR_253 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_3_NAND3X1_25 DFFSR_8/gnd DFFSR_8/S FILL
XDFFSR_143 DFFSR_143/Q CLKBUF1_20/Y BUFX2_62/Y DFFSR_216/S DFFSR_183/Q OR2X2_2/gnd
+ DFFSR_216/S DFFSR
XFILL_2_NAND3X1_28 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_3_OAI22X1_10 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_29_6_1 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_14_DFFSR_35 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_4_DFFSR_140 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_1_BUFX2_70 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_1_NAND3X1_31 BUFX2_79/A DFFSR_6/S FILL
XFILL_2_OAI22X1_13 INVX1_1/gnd DFFSR_53/S FILL
XFILL_45_DFFSR_171 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_0_NAND3X1_34 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_8_DFFSR_247 BUFX2_99/A DFFSR_7/S FILL
XFILL_1_OAI22X1_16 AND2X2_38/B DFFSR_59/S FILL
XFILL_35_DFFSR_174 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_23_DFFPOSX1_10 INVX1_67/gnd DFFSR_201/S FILL
XFILL_49_DFFSR_278 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_0_OAI22X1_19 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_45_DFFSR_2 BUFX2_79/A DFFSR_7/S FILL
XFILL_25_DFFSR_177 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_49_DFFSR_52 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_38_DFFSR_92 BUFX2_99/A DFFSR_92/S FILL
XFILL_15_DFFSR_180 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_7_NAND3X1_213 INVX1_39/gnd DFFSR_54/S FILL
XFILL_3_DFFPOSX1_32 INVX1_67/gnd DFFSR_201/S FILL
XINVX1_36 INVX1_36/A OR2X2_3/gnd INVX1_36/Y DFFSR_4/S INVX1
XDFFSR_89 DFFSR_89/Q CLKBUF1_18/Y DFFSR_73/R DFFSR_59/S INVX1_5/A OR2X2_1/gnd DFFSR_59/S
+ DFFSR
XFILL_22_DFFSR_42 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_5_DFFSR_49 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_11_DFFSR_82 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_0_NOR2X1_59 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_2_OAI21X1_7 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_38_DFFSR_101 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_8_NAND3X1_147 OR2X2_1/gnd DFFSR_51/S FILL
XINVX1_154 INVX1_154/A XOR2X1_1/gnd INVX1_154/Y DFFSR_208/S INVX1
XFILL_0_INVX1_4 BUFX2_99/A DFFSR_7/S FILL
XFILL_1_6 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_1_DFFSR_177 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_28_DFFSR_104 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_1_NAND2X1_128 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_42_DFFSR_208 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_46_DFFSR_99 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_7_AND2X2_18 AND2X2_38/B DFFSR_59/S FILL
XFILL_18_DFFSR_107 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_32_DFFSR_211 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_22_DFFSR_214 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_7_AND2X2_8 BUFX2_99/A DFFSR_7/S FILL
XFILL_2_INVX1_43 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_2_DFFSR_96 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_30_DFFSR_49 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_19_DFFSR_89 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_39_1_1 BUFX2_79/A DFFSR_6/S FILL
XFILL_12_DFFSR_217 BUFX2_72/gnd DFFSR_201/S FILL
XDFFSR_107 DFFSR_115/D DFFSR_9/CLK DFFSR_73/R DFFSR_92/S DFFSR_99/Q OR2X2_6/gnd DFFSR_92/S
+ DFFSR
XFILL_22_DFFPOSX1_40 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_4_DFFSR_104 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_37_3_2 BUFX2_99/A DFFSR_7/S FILL
XFILL_6_NAND3X1_243 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_1_BUFX2_34 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_45_DFFSR_135 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_8_DFFSR_211 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_35_DFFSR_138 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_49_DFFSR_242 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_25_DFFSR_141 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_39_DFFSR_245 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_49_DFFSR_16 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_38_DFFSR_56 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_27_DFFSR_96 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_1_INVX1_188 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_1_CLKBUF1_9 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_7_NAND3X1_177 AND2X2_38/B DFFSR_59/S FILL
XFILL_15_DFFSR_144 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_29_DFFSR_248 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_19_DFFSR_251 BUFX2_7/gnd DFFSR_151/S FILL
XDFFSR_53 INVX1_31/A DFFSR_9/CLK BUFX2_49/Y DFFSR_53/S INVX1_32/A OR2X2_6/gnd DFFSR_53/S
+ DFFSR
XFILL_0_NAND2X1_158 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_5_DFFSR_13 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_11_DFFSR_46 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_0_NOR2X1_23 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_8_NAND3X1_111 XOR2X1_1/gnd DFFSR_151/S FILL
XINVX1_118 BUFX2_40/Y BUFX2_98/A BUFX2_60/A DFFSR_6/S INVX1
XFILL_12_DFFPOSX1_15 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_1_DFFSR_141 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_4_INVX1_115 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_42_DFFSR_172 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_46_DFFSR_63 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_5_DFFSR_248 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_32_DFFSR_175 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_46_DFFSR_279 BUFX2_99/A DFFSR_7/S FILL
XFILL_22_DFFSR_178 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_2_DFFSR_60 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_30_DFFSR_13 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_19_DFFSR_53 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_12_DFFSR_181 INVX1_3/gnd DFFSR_79/S FILL
XFILL_6_BUFX2_88 INVX1_3/gnd DFFSR_23/S FILL
XFILL_20_CLKBUF1_43 AND2X2_38/B DFFSR_23/S FILL
XFILL_6_NAND3X1_207 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_19_CLKBUF1_46 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_36_DFFSR_9 BUFX2_79/A DFFSR_6/S FILL
XFILL_2_DFFPOSX1_26 AND2X2_38/B DFFSR_23/S FILL
XFILL_8_DFFSR_175 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_35_DFFSR_102 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_49_DFFSR_206 OR2X2_2/gnd DFFSR_175/S FILL
XAND2X2_22 AND2X2_22/A AND2X2_22/B OR2X2_1/gnd AND2X2_22/Y DFFSR_59/S AND2X2
XFILL_18_CLKBUF1_49 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_25_DFFSR_105 INVX1_1/gnd DFFSR_53/S FILL
XNAND3X1_243 XOR2X1_8/A NAND3X1_243/B NAND3X1_242/Y DFFSR_28/gnd AOI21X1_45/B DFFSR_3/S
+ NAND3X1
XFILL_39_DFFSR_209 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_27_DFFSR_60 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_38_DFFSR_20 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_1_INVX1_152 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_4_AND2X2_19 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_15_DFFSR_108 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_7_NAND3X1_141 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_29_DFFSR_212 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_11_DFFPOSX1_45 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_0_NAND2X1_122 INVX1_67/gnd DFFSR_175/S FILL
XDFFSR_17 INVX1_7/A CLKBUF1_7/Y DFFSR_3/R DFFSR_3/S INVX1_8/A DFFSR_28/gnd DFFSR_3/S
+ DFFSR
XFILL_19_DFFSR_215 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_11_DFFSR_10 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_1_DFFSR_105 INVX1_1/gnd DFFSR_53/S FILL
XFILL_21_DFFPOSX1_34 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_42_DFFSR_136 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_11_1_2 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_46_DFFSR_27 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_35_DFFSR_67 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_5_DFFSR_212 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_32_DFFSR_139 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_46_DFFSR_243 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_5_NAND3X1_237 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_8_CLKBUF1_7 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_22_DFFSR_142 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_2_DFFSR_24 BUFX2_98/A DFFSR_6/S FILL
XFILL_36_DFFSR_246 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_19_DFFSR_17 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_12_DFFSR_145 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_6_BUFX2_52 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_26_DFFSR_249 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_16_DFFSR_252 AND2X2_38/B DFFSR_23/S FILL
XFILL_1_NOR2X1_5 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_6_NAND3X1_171 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_19_CLKBUF1_10 INVX1_67/gnd DFFSR_201/S FILL
XFILL_43_DFFSR_74 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_8_DFFSR_139 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_18_CLKBUF1_13 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_49_DFFSR_170 OR2X2_6/gnd DFFSR_92/S FILL
XNAND3X1_207 INVX1_164/A OAI21X1_71/Y OAI21X1_72/Y DFFSR_1/gnd NAND3X1_214/A DFFSR_1/S
+ NAND3X1
XFILL_17_CLKBUF1_16 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_39_DFFSR_173 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_1_INVX1_116 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_27_DFFSR_24 BUFX2_98/A DFFSR_6/S FILL
XFILL_16_DFFSR_64 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_38_4_0 BUFX2_79/A DFFSR_7/S FILL
XFILL_2_DFFSR_249 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_7_NAND3X1_105 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_3_BUFX2_99 BUFX2_99/A DFFSR_7/S FILL
XFILL_29_DFFSR_176 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_16_CLKBUF1_19 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_43_DFFSR_280 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_15_CLKBUF1_22 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_19_DFFSR_179 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_36_6_1 BUFX2_99/A DFFSR_92/S FILL
XNOR2X1_61 NOR3X1_4/B NOR3X1_4/A BUFX2_8/gnd NOR2X1_61/Y DFFSR_51/S NOR2X1
XFILL_14_CLKBUF1_25 INVX1_67/gnd DFFSR_201/S FILL
XFILL_3_XOR2X1_1 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_13_CLKBUF1_28 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_23_DFFSR_3 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_51_DFFSR_81 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_4_NOR2X1_58 INVX1_3/gnd DFFSR_79/S FILL
XFILL_6_OAI21X1_6 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_12_CLKBUF1_31 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_42_DFFSR_100 INVX1_1/gnd DFFSR_97/S FILL
XFILL_7_DFFSR_78 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_11_CLKBUF1_34 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_35_DFFSR_31 BUFX2_79/A DFFSR_6/S FILL
XFILL_24_DFFSR_71 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_5_DFFSR_176 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_32_DFFSR_103 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_10_CLKBUF1_37 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_5_NAND3X1_201 INVX1_1/gnd DFFSR_53/S FILL
XFILL_46_DFFSR_207 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_22_DFFSR_106 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_36_DFFSR_210 BUFX2_98/A DFFSR_6/S FILL
XFILL_1_DFFPOSX1_20 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_1_AND2X2_20 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_12_DFFSR_109 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_6_BUFX2_16 BUFX2_98/A DFFSR_32/S FILL
XFILL_9_CLKBUF1_40 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_26_DFFSR_213 INVX1_3/gnd DFFSR_23/S FILL
XFILL_16_DFFSR_216 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_8_CLKBUF1_43 AND2X2_38/B DFFSR_23/S FILL
XFILL_6_NAND3X1_135 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_7_CLKBUF1_46 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_10_DFFPOSX1_39 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_32_DFFSR_78 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_43_DFFSR_38 BUFX2_98/A DFFSR_6/S FILL
XFILL_4_INVX1_72 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_8_DFFSR_103 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_6_CLKBUF1_49 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_49_DFFSR_134 INVX1_1/gnd DFFSR_53/S FILL
XNAND3X1_171 OAI21X1_47/Y INVX1_158/Y NAND2X1_83/Y DFFSR_34/gnd AOI22X1_23/A DFFSR_34/S
+ NAND3X1
XFILL_39_DFFSR_137 BUFX2_7/gnd DFFSR_216/S FILL
XCLKBUF1_49 clk BUFX2_8/gnd CLKBUF1_49/Y DFFSR_81/S CLKBUF1
XFILL_16_DFFSR_28 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_2_DFFSR_213 INVX1_3/gnd DFFSR_23/S FILL
XFILL_3_BUFX2_63 BUFX2_98/A DFFSR_32/S FILL
XFILL_29_DFFSR_140 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_46_1_1 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_43_DFFSR_244 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_20_DFFPOSX1_28 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_19_DFFSR_143 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_5_CLKBUF1_8 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_33_DFFSR_247 BUFX2_99/A DFFSR_7/S FILL
XNOR2X1_25 NOR2X1_25/A NOR2X1_25/B DFFSR_28/gnd NOR2X1_25/Y DFFSR_8/S NOR2X1
XFILL_44_3_2 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_23_DFFSR_250 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_4_NAND3X1_231 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_51_DFFSR_45 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_40_DFFSR_85 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_4_NOR2X1_22 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_0_DFFPOSX1_50 INVX1_1/gnd DFFSR_53/S FILL
XFILL_13_DFFSR_253 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_7_DFFSR_42 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_24_DFFSR_35 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_13_DFFSR_75 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_5_DFFSR_140 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_46_DFFSR_171 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_5_NAND3X1_165 INVX1_39/gnd DFFSR_34/S FILL
XFILL_9_DFFSR_247 BUFX2_99/A DFFSR_7/S FILL
XFILL_36_DFFSR_174 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_50_DFFSR_278 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_26_DFFSR_177 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_12_2_0 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_48_DFFSR_92 BUFX2_99/A DFFSR_92/S FILL
XFILL_16_DFFSR_180 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_7_CLKBUF1_10 INVX1_67/gnd DFFSR_201/S FILL
XFILL_9_AND2X2_1 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_10_4_1 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_4_INVX1_36 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_32_DFFSR_42 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_4_DFFSR_89 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_21_DFFSR_82 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_6_CLKBUF1_13 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_1_NOR2X1_59 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_3_OAI21X1_7 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_5_CLKBUF1_16 OR2X2_3/gnd DFFSR_4/S FILL
XNAND3X1_135 BUFX2_7/Y OR2X2_1/A NOR3X1_1/A BUFX2_8/gnd NAND2X1_57/B DFFSR_81/S NAND3X1
XFILL_39_DFFSR_101 OR2X2_3/gnd DFFSR_4/S FILL
XCLKBUF1_13 BUFX2_1/Y DFFSR_28/gnd DFFSR_8/CLK DFFSR_3/S CLKBUF1
XFILL_5_3 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_4_CLKBUF1_19 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_2_DFFSR_177 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_29_DFFSR_104 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_3_BUFX2_27 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_43_DFFSR_208 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_3_CLKBUF1_22 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_8_AND2X2_18 AND2X2_38/B DFFSR_59/S FILL
XFILL_19_DFFSR_107 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_6_OAI21X1_117 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_2_CLKBUF1_25 INVX1_67/gnd DFFSR_201/S FILL
XFILL_33_DFFSR_211 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_13_NOR3X1_6 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_23_DFFSR_214 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_1_CLKBUF1_28 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_4_NAND3X1_195 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_40_DFFSR_49 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_29_DFFSR_89 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_1_INVX1_83 INVX1_39/gnd DFFSR_54/S FILL
XFILL_13_DFFSR_217 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_0_CLKBUF1_31 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_0_DFFPOSX1_14 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_13_DFFSR_39 INVX1_3/gnd DFFSR_79/S FILL
XFILL_5_DFFSR_104 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_0_BUFX2_74 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_9_OR2X2_2 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_5_NAND3X1_129 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_46_DFFSR_135 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_9_DFFSR_211 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_36_DFFSR_138 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_50_DFFSR_242 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_35_DFFSR_6 BUFX2_79/A DFFSR_6/S FILL
XFILL_26_DFFSR_141 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_40_DFFSR_245 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_48_DFFSR_56 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_37_DFFSR_96 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_2_INVX1_188 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_2_CLKBUF1_9 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_16_DFFSR_144 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_30_DFFSR_248 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_20_DFFSR_251 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_4_DFFSR_53 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_10_DFFSR_86 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_19_DFFPOSX1_22 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_18_1_2 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_21_DFFSR_46 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_1_NOR2X1_23 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_10_DFFSR_254 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_0_0_1 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_3_NAND3X1_225 DFFSR_4/gnd DFFSR_4/S FILL
XBUFX2_100 BUFX2_79/A BUFX2_79/A BUFX2_100/Y DFFSR_6/S BUFX2
XFILL_2_DFFSR_141 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_43_DFFSR_172 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_6_DFFSR_248 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_33_DFFSR_175 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_47_DFFSR_279 BUFX2_99/A DFFSR_7/S FILL
XFILL_23_DFFSR_178 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_4_NAND3X1_159 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_18_DFFSR_93 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_1_INVX1_47 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_40_DFFSR_13 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_29_DFFSR_53 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_13_DFFSR_181 INVX1_3/gnd DFFSR_79/S FILL
XOAI21X1_117 XOR2X1_14/Y OAI21X1_116/Y AOI21X1_69/Y XOR2X1_4/gnd NOR2X1_82/B DFFSR_97/S
+ OAI21X1
XFILL_9_DFFPOSX1_33 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_0_BUFX2_38 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_45_4_0 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_0_OAI21X1_8 BUFX2_99/A DFFSR_7/S FILL
XFILL_9_DFFSR_175 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_36_DFFSR_102 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_50_DFFSR_206 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_43_6_1 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_26_DFFSR_105 INVX1_1/gnd DFFSR_53/S FILL
XFILL_40_DFFSR_209 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_37_DFFSR_60 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_48_DFFSR_20 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_2_INVX1_152 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_5_AND2X2_19 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_16_DFFSR_108 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_30_DFFSR_212 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_20_DFFSR_215 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_4_DFFSR_17 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_21_DFFSR_10 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_10_DFFSR_50 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_5_OAI21X1_111 AND2X2_38/B DFFSR_59/S FILL
XFILL_10_DFFSR_218 BUFX2_98/A DFFSR_32/S FILL
XFILL_3_NAND3X1_189 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_2_DFFSR_9 BUFX2_79/A DFFSR_6/S FILL
XFILL_2_DFFSR_105 INVX1_1/gnd DFFSR_53/S FILL
XFILL_43_DFFSR_136 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_45_DFFSR_67 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_6_DFFSR_212 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_33_DFFSR_139 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_47_DFFSR_243 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_23_DFFSR_142 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_9_CLKBUF1_7 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_4_NAND3X1_123 BUFX2_99/A DFFSR_7/S FILL
XFILL_29_DFFSR_17 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_1_DFFSR_64 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_1_INVX1_11 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_18_DFFSR_57 BUFX2_79/A DFFSR_6/S FILL
XFILL_37_DFFSR_246 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_13_DFFSR_145 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_5_BUFX2_92 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_6_BUFX2_1 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_27_DFFSR_249 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_6_NAND2X1_159 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_49_4 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_17_DFFSR_252 AND2X2_38/B DFFSR_23/S FILL
XFILL_53_1_1 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_9_DFFSR_139 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_18_DFFPOSX1_16 INVX1_67/gnd DFFSR_175/S FILL
XFILL_50_DFFSR_170 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_40_DFFSR_173 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_51_3_2 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_2_INVX1_116 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_37_DFFSR_24 BUFX2_98/A DFFSR_6/S FILL
XFILL_9_DFFSR_71 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_26_DFFSR_64 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_3_DFFSR_249 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_18_DFFPOSX1_1 INVX1_39/gnd DFFSR_34/S FILL
XFILL_2_NAND3X1_219 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_30_DFFSR_176 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_44_DFFSR_280 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_17_DFFPOSX1_4 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_20_DFFSR_179 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_10_DFFSR_14 INVX1_1/gnd DFFSR_53/S FILL
XFILL_16_DFFPOSX1_7 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_10_DFFSR_182 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_5_NOR2X1_58 INVX1_3/gnd DFFSR_79/S FILL
XFILL_3_NAND3X1_153 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_47_DFFSR_9 BUFX2_79/A DFFSR_6/S FILL
XFILL_7_OAI21X1_6 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_43_DFFSR_100 INVX1_1/gnd DFFSR_97/S FILL
XFILL_8_DFFPOSX1_27 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_45_DFFSR_31 BUFX2_79/A DFFSR_6/S FILL
XFILL_34_DFFSR_71 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_19_2_0 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_6_DFFSR_176 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_33_DFFSR_103 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_47_DFFSR_207 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_23_DFFSR_106 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_1_DFFSR_28 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_18_DFFSR_21 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_37_DFFSR_210 BUFX2_98/A DFFSR_6/S FILL
XFILL_17_4_1 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_2_AND2X2_20 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_13_DFFSR_109 DFFSR_4/gnd DFFSR_4/S FILL
XBUFX2_96 BUFX2_96/A OR2X2_4/gnd BUFX2_96/Y DFFSR_32/S BUFX2
XFILL_5_BUFX2_56 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_17_DFFPOSX1_46 INVX1_39/gnd DFFSR_34/S FILL
XFILL_10_OAI22X1_2 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_27_DFFSR_213 INVX1_3/gnd DFFSR_23/S FILL
XFILL_6_NAND2X1_123 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_17_DFFSR_216 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_9_NOR3X1_2 INVX1_1/gnd DFFSR_53/S FILL
XFILL_0_NOR2X1_9 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_1_NAND3X1_249 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_15_6_2 INVX1_39/gnd DFFSR_34/S FILL
XFILL_9_DFFSR_103 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_42_DFFSR_78 OR2X2_3/gnd DFFSR_4/S FILL
XNAND2X1_159 DFFSR_91/S NAND2X1_160/A XOR2X1_4/gnd AOI21X1_55/B DFFSR_91/S NAND2X1
XFILL_4_OAI21X1_105 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_50_DFFSR_134 INVX1_1/gnd DFFSR_53/S FILL
XFILL_8_AOI21X1_51 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_27_DFFPOSX1_35 INVX1_39/gnd DFFSR_54/S FILL
XFILL_40_DFFSR_137 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_9_DFFSR_35 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_7_AOI21X1_54 AND2X2_38/B DFFSR_59/S FILL
XFILL_26_DFFSR_28 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_15_DFFSR_68 BUFX2_98/A DFFSR_6/S FILL
XFILL_3_DFFSR_213 INVX1_3/gnd DFFSR_23/S FILL
XFILL_2_NAND3X1_183 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_30_DFFSR_140 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_6_AOI21X1_57 INVX1_67/gnd DFFSR_201/S FILL
XFILL_44_DFFSR_244 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_20_DFFSR_143 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_6_CLKBUF1_8 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_5_AOI21X1_60 BUFX2_79/A DFFSR_7/S FILL
XFILL_34_DFFSR_247 BUFX2_99/A DFFSR_7/S FILL
XAOI21X1_57 AOI21X1_57/A AOI21X1_57/B BUFX2_36/Y INVX1_67/gnd AOI21X1_57/Y DFFSR_201/S
+ AOI21X1
XFILL_10_DFFSR_146 BUFX2_79/A DFFSR_7/S FILL
XFILL_4_AOI21X1_63 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_24_DFFSR_250 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_2_XOR2X1_5 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_50_DFFSR_85 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_5_NOR2X1_22 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_13_DFFSR_7 BUFX2_79/A DFFSR_7/S FILL
XFILL_3_NAND3X1_117 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_3_AOI21X1_66 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_14_DFFSR_253 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_2_AOI21X1_69 INVX1_1/gnd DFFSR_97/S FILL
XFILL_34_DFFSR_35 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_6_DFFSR_82 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_5_NAND2X1_153 BUFX2_98/A DFFSR_32/S FILL
XFILL_23_DFFSR_75 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_6_DFFSR_140 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_47_DFFSR_171 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_37_DFFSR_174 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_51_DFFSR_278 XOR2X1_1/gnd DFFSR_151/S FILL
XBUFX2_60 BUFX2_60/A OR2X2_2/gnd BUFX2_60/Y DFFSR_216/S BUFX2
XFILL_0_DFFSR_250 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_5_BUFX2_20 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_17_DFFPOSX1_10 INVX1_67/gnd DFFSR_201/S FILL
XFILL_25_1_2 AND2X2_38/B DFFSR_23/S FILL
XFILL_27_DFFSR_177 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_9_OAI21X1_96 AND2X2_38/B DFFSR_59/S FILL
XFILL_17_DFFSR_180 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_7_0_1 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_8_OAI21X1_99 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_34_DFFSR_3 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_1_NAND3X1_213 INVX1_39/gnd DFFSR_54/S FILL
XFILL_42_DFFSR_42 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_3_INVX1_76 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_31_DFFSR_82 BUFX2_77/gnd DFFSR_98/S FILL
XNAND2X1_123 DFFSR_264/S din[7] BUFX2_77/gnd OAI21X1_92/C DFFSR_98/S NAND2X1
XFILL_2_NOR2X1_59 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_5_2_2 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_4_OAI21X1_7 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_8_AOI21X1_15 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_40_DFFSR_101 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_7_AOI21X1_18 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_6_DFFPOSX1_1 INVX1_39/gnd DFFSR_34/S FILL
XFILL_15_DFFSR_32 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_2_NAND3X1_147 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_3_DFFSR_177 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_2_BUFX2_67 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_30_DFFSR_104 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_5_DFFPOSX1_4 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_6_AOI21X1_21 INVX1_39/gnd DFFSR_54/S FILL
XFILL_44_DFFSR_208 DFFSR_62/gnd DFFSR_208/S FILL
XDFFPOSX1_1 BUFX2_3/A CLKBUF1_49/Y DFFPOSX1_1/D INVX1_39/gnd DFFSR_34/S DFFPOSX1
XFILL_7_DFFPOSX1_21 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_20_DFFSR_107 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_4_DFFPOSX1_7 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_5_AOI21X1_24 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_34_DFFSR_211 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_10_DFFSR_110 OR2X2_3/gnd DFFSR_4/S FILL
XAOI21X1_21 AOI21X1_21/A AOI21X1_21/B OAI21X1_58/C INVX1_39/gnd OAI21X1_54/B DFFSR_54/S
+ AOI21X1
XFILL_4_AOI21X1_27 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_24_DFFSR_214 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_52_4_0 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_50_DFFSR_49 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_39_DFFSR_89 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_14_DFFSR_217 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_3_AOI21X1_30 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_16_DFFPOSX1_40 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_2_AOI21X1_33 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_50_6_1 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_5_NAND2X1_117 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_23_DFFSR_39 INVX1_3/gnd DFFSR_79/S FILL
XFILL_6_DFFSR_46 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_6_DFFSR_104 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_1_AOI21X1_36 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_12_DFFSR_79 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_0_NAND3X1_243 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_47_DFFSR_135 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_0_AOI21X1_39 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_37_DFFSR_138 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_51_DFFSR_242 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_0_DFFSR_214 BUFX2_72/gnd DFFSR_276/S FILL
XBUFX2_24 BUFX2_23/A XOR2X1_1/gnd BUFX2_24/Y DFFSR_151/S BUFX2
XFILL_27_DFFSR_141 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_26_DFFPOSX1_29 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_31_1 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_3_INVX1_188 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_41_DFFSR_245 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_47_DFFSR_96 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_3_CLKBUF1_9 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_17_DFFSR_144 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_8_OAI21X1_63 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_31_DFFSR_248 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_1_NAND3X1_177 AND2X2_38/B DFFSR_59/S FILL
XFILL_21_DFFSR_251 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_8_AND2X2_5 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_7_OAI21X1_66 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_6_NAND2X1_84 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_3_INVX1_40 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_3_DFFSR_93 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_20_DFFSR_86 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_31_DFFSR_46 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_2_NOR2X1_23 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_5_NAND2X1_87 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_6_OAI21X1_69 INVX1_3/gnd DFFSR_23/S FILL
XFILL_11_DFFSR_254 DFFSR_34/gnd DFFSR_1/S FILL
XNAND2X1_84 INVX1_175/A AND2X2_34/B NOR3X1_6/gnd INVX1_160/A DFFSR_91/S NAND2X1
XFILL_5_OAI21X1_72 INVX1_3/gnd DFFSR_23/S FILL
XFILL_4_NAND2X1_90 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_2_NAND3X1_111 XOR2X1_1/gnd DFFSR_151/S FILL
XOAI21X1_69 OAI21X1_69/A OAI21X1_69/B OAI21X1_61/Y INVX1_3/gnd OAI21X1_69/Y DFFSR_23/S
+ OAI21X1
XFILL_3_NAND2X1_93 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_3_DFFSR_141 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_4_OAI21X1_75 INVX1_39/gnd DFFSR_54/S FILL
XFILL_2_BUFX2_31 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_44_DFFSR_172 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_3_OAI21X1_78 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_2_NAND2X1_96 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_7_DFFSR_248 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_1_DFFSR_6 BUFX2_79/A DFFSR_6/S FILL
XFILL_4_NAND2X1_147 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_34_DFFSR_175 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_2_OAI21X1_81 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_1_NAND2X1_99 INVX1_39/gnd DFFSR_54/S FILL
XFILL_48_DFFSR_279 BUFX2_99/A DFFSR_7/S FILL
XFILL_24_DFFSR_178 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_1_OAI21X1_84 BUFX2_98/A DFFSR_6/S FILL
XFILL_0_INVX1_87 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_50_DFFSR_13 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_39_DFFSR_53 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_28_DFFSR_93 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_14_DFFSR_181 INVX1_3/gnd DFFSR_79/S FILL
XFILL_0_OAI21X1_87 BUFX2_79/A DFFSR_7/S FILL
XFILL_6_DFFSR_10 DFFSR_5/gnd DFFSR_5/S FILL
XBUFX2_2 BUFX2_3/A OR2X2_4/gnd BUFX2_2/Y DFFSR_32/S BUFX2
XFILL_12_DFFSR_43 BUFX2_98/A DFFSR_6/S FILL
XFILL_1_OAI21X1_8 BUFX2_99/A DFFSR_7/S FILL
XFILL_0_NAND3X1_207 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_37_DFFSR_102 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_0_DFFSR_178 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_27_DFFSR_105 INVX1_1/gnd DFFSR_53/S FILL
XFILL_9_OAI21X1_24 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_41_DFFSR_209 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_3_INVX1_152 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_6_AND2X2_19 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_47_DFFSR_60 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_17_DFFSR_108 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_8_OAI21X1_27 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_31_DFFSR_212 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_1_NAND3X1_141 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_6_NAND2X1_48 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_7_OAI21X1_30 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_21_DFFSR_215 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_3_DFFSR_57 BUFX2_79/A DFFSR_6/S FILL
XFILL_31_DFFSR_10 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_20_DFFSR_50 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_6_DFFPOSX1_15 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_11_DFFSR_218 BUFX2_98/A DFFSR_32/S FILL
XFILL_3_NAND2X1_177 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_5_NAND2X1_51 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_6_OAI21X1_33 INVX1_3/gnd DFFSR_79/S FILL
XFILL_26_2_0 INVX1_3/gnd DFFSR_23/S FILL
XNAND2X1_48 DFFSR_174/D AND2X2_18/Y BUFX2_8/gnd NAND2X1_48/Y DFFSR_81/S NAND2X1
XFILL_4_NAND2X1_54 AND2X2_38/B DFFSR_59/S FILL
XFILL_5_OAI21X1_36 BUFX2_8/gnd DFFSR_51/S FILL
XOAI21X1_33 INVX1_132/Y INVX1_146/Y AND2X2_31/Y INVX1_3/gnd OAI21X1_33/Y DFFSR_79/S
+ OAI21X1
XFILL_3_DFFSR_105 INVX1_1/gnd DFFSR_53/S FILL
XFILL_3_NAND2X1_57 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_4_OAI21X1_39 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_24_4_1 AND2X2_38/B DFFSR_59/S FILL
XFILL_44_DFFSR_136 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_15_DFFPOSX1_34 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_3_OAI21X1_42 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_46_DFFSR_6 BUFX2_79/A DFFSR_6/S FILL
XFILL_2_NAND2X1_60 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_7_DFFSR_212 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_6_3_0 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_4_NAND2X1_111 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_34_DFFSR_139 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_48_DFFSR_243 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_1_NAND2X1_63 AND2X2_38/B DFFSR_59/S FILL
XFILL_2_OAI21X1_45 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_11_AOI22X1_11 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_22_6_2 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_24_DFFSR_142 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_1_OAI21X1_48 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_0_NAND2X1_66 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_10_AOI22X1_14 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_39_DFFSR_17 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_0_INVX1_51 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_28_DFFSR_57 BUFX2_79/A DFFSR_6/S FILL
XFILL_0_INVX1_189 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_38_DFFSR_246 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_17_DFFSR_97 INVX1_1/gnd DFFSR_97/S FILL
XFILL_14_DFFSR_145 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_4_5_1 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_0_OAI21X1_51 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_28_DFFSR_249 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_36_6 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_53_1 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_25_DFFPOSX1_23 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_18_DFFSR_252 AND2X2_38/B DFFSR_23/S FILL
XFILL_9_AOI22X1_17 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_1_INVX1_8 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_0_NAND3X1_171 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_8_AOI22X1_20 INVX1_39/gnd DFFSR_34/S FILL
XFILL_7_AOI22X1_23 INVX1_39/gnd DFFSR_34/S FILL
XFILL_51_DFFSR_170 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_5_DFFPOSX1_45 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_0_DFFSR_142 XOR2X1_1/gnd DFFSR_151/S FILL
XDFFSR_252 BUFX2_93/A CLKBUF1_18/Y BUFX2_61/Y DFFSR_23/S INVX1_89/A AND2X2_38/B DFFSR_23/S
+ DFFSR
XFILL_6_AOI22X1_26 INVX1_1/gnd DFFSR_97/S FILL
XFILL_3_INVX1_116 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_41_DFFSR_173 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_36_DFFSR_64 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_47_DFFSR_24 BUFX2_98/A DFFSR_6/S FILL
XFILL_4_DFFSR_249 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_5_AOI22X1_29 INVX1_1/gnd DFFSR_53/S FILL
XFILL_31_DFFSR_176 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_1_NAND3X1_105 DFFSR_1/gnd DFFSR_81/S FILL
XAOI22X1_26 AOI22X1_26/A AOI22X1_26/B AOI22X1_26/C AOI22X1_26/D INVX1_1/gnd OAI21X1_69/A
+ DFFSR_97/S AOI22X1
XFILL_45_DFFSR_280 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_6_NAND2X1_12 INVX1_3/gnd DFFSR_79/S FILL
XFILL_21_DFFSR_179 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_3_DFFSR_21 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_20_DFFSR_14 INVX1_1/gnd DFFSR_53/S FILL
XFILL_5_NAND2X1_15 BUFX2_99/A DFFSR_92/S FILL
XFILL_3_NAND2X1_141 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_11_DFFSR_182 XOR2X1_1/gnd DFFSR_208/S FILL
XNAND2X1_12 OR2X2_1/A BUFX2_8/Y INVX1_3/gnd NOR3X1_1/C DFFSR_79/S NAND2X1
XFILL_4_NAND2X1_18 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_6_NOR2X1_58 INVX1_3/gnd DFFSR_79/S FILL
XFILL_8_OAI21X1_6 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_3_NAND2X1_21 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_2_NOR2X1_2 INVX1_1/gnd DFFSR_97/S FILL
XDFFPOSX1_15 INVX1_137/A CLKBUF1_47/Y OAI21X1_23/Y BUFX2_72/gnd DFFSR_201/S DFFPOSX1
XFILL_12_DFFSR_4 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_44_DFFSR_100 INVX1_1/gnd DFFSR_97/S FILL
XFILL_2_NAND2X1_24 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_32_1_2 INVX1_1/gnd DFFSR_97/S FILL
XFILL_44_DFFSR_71 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_7_DFFSR_176 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_34_DFFSR_103 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_1_NAND2X1_27 AND2X2_38/B DFFSR_23/S FILL
XFILL_48_DFFSR_207 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_8_NAND3X1_83 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_24_DFFSR_106 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_0_NAND2X1_30 AND2X2_38/B DFFSR_23/S FILL
XFILL_1_OAI21X1_12 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_0_INVX1_153 INVX1_67/gnd DFFSR_175/S FILL
XFILL_28_DFFSR_21 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_0_INVX1_15 BUFX2_98/A DFFSR_32/S FILL
XFILL_0_DFFSR_68 BUFX2_98/A DFFSR_6/S FILL
XFILL_38_DFFSR_210 BUFX2_98/A DFFSR_6/S FILL
XFILL_17_DFFSR_61 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_3_AND2X2_20 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_14_DFFSR_109 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_7_NAND3X1_86 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_4_BUFX2_96 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_0_OAI21X1_15 INVX1_3/gnd DFFSR_79/S FILL
XFILL_28_DFFSR_213 INVX1_3/gnd DFFSR_23/S FILL
XFILL_6_NAND3X1_89 DFFSR_62/gnd DFFSR_62/S FILL
XFILL_18_DFFSR_216 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_5_NAND3X1_92 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_0_NAND3X1_135 BUFX2_8/gnd DFFSR_81/S FILL
XNAND3X1_89 DFFSR_172/Q BUFX2_27/Y BUFX2_23/Y DFFSR_62/gnd NAND3X1_89/Y DFFSR_62/S
+ NAND3X1
XFILL_4_NAND3X1_95 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_51_DFFSR_134 INVX1_1/gnd DFFSR_53/S FILL
XDFFSR_216 DFFSR_216/Q CLKBUF1_10/Y BUFX2_64/Y DFFSR_216/S DFFSR_216/D BUFX2_7/gnd
+ DFFSR_216/S DFFSR
XFILL_0_DFFSR_106 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_3_NAND3X1_98 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_2_NAND2X1_171 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_41_DFFSR_137 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_36_DFFSR_28 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_25_DFFSR_68 BUFX2_98/A DFFSR_6/S FILL
XFILL_8_DFFSR_75 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_4_DFFSR_213 INVX1_3/gnd DFFSR_23/S FILL
XFILL_31_DFFSR_140 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_45_DFFSR_244 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_21_DFFSR_143 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_7_CLKBUF1_8 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_14_DFFPOSX1_28 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_35_DFFSR_247 BUFX2_99/A DFFSR_7/S FILL
XFILL_11_DFFSR_146 BUFX2_79/A DFFSR_7/S FILL
XFILL_3_NAND2X1_105 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_25_DFFSR_250 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_6_NOR2X1_22 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_15_DFFSR_253 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_10_OAI22X1_26 INVX1_39/gnd DFFSR_54/S FILL
XFILL_44_DFFSR_35 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_33_DFFSR_75 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_7_DFFSR_140 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_24_DFFPOSX1_17 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_9_NAND3X1_44 BUFX2_99/A DFFSR_7/S FILL
XFILL_48_DFFSR_171 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_8_NAND3X1_47 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_9_OAI22X1_29 INVX1_3/gnd DFFSR_79/S FILL
XFILL_0_INVX1_117 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_0_DFFSR_32 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_38_DFFSR_174 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_8_NAND3X1_220 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_17_DFFSR_25 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_1_DFFSR_250 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_7_NAND3X1_50 BUFX2_98/A DFFSR_6/S FILL
XFILL_8_OAI22X1_32 INVX1_39/gnd DFFSR_54/S FILL
XFILL_4_BUFX2_60 OR2X2_2/gnd DFFSR_216/S FILL
XFILL_4_DFFPOSX1_39 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_28_DFFSR_177 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_6_NAND3X1_53 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_7_OAI22X1_35 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_18_DFFSR_180 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_8_NOR3X1_6 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_5_NAND3X1_56 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_6_OAI22X1_38 AND2X2_38/B DFFSR_23/S FILL
XNAND3X1_53 DFFSR_71/D BUFX2_19/Y BUFX2_13/Y OR2X2_3/gnd NAND3X1_53/Y DFFSR_60/S NAND3X1
XFILL_9_NAND3X1_154 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_4_NAND3X1_59 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_5_OAI22X1_41 INVX1_39/gnd DFFSR_54/S FILL
XFILL_41_DFFSR_82 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_3_NOR2X1_59 DFFSR_34/gnd DFFSR_1/S FILL
XOAI22X1_38 INVX1_92/Y OAI22X1_41/B INVX1_93/Y OAI22X1_41/D AND2X2_38/B NOR2X1_47/A
+ DFFSR_23/S OAI22X1
XFILL_5_OAI21X1_7 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_3_NAND3X1_62 DFFSR_8/gnd DFFSR_60/S FILL
XFILL_4_OAI22X1_44 DFFSR_1/gnd DFFSR_81/S FILL
XDFFSR_180 INVX1_83/A DFFSR_1/CLK BUFX2_69/Y DFFSR_34/S INVX1_84/A DFFSR_34/gnd DFFSR_34/S
+ DFFSR
XFILL_2_NAND2X1_135 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_41_DFFSR_101 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_3_OAI22X1_47 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_2_NAND3X1_65 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_14_DFFSR_72 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_25_DFFSR_32 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_8_DFFSR_39 INVX1_3/gnd DFFSR_79/S FILL
XFILL_4_DFFSR_177 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_1_NAND3X1_68 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_31_DFFSR_104 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_2_OAI22X1_50 INVX1_3/gnd DFFSR_23/S FILL
XFILL_45_DFFSR_208 DFFSR_62/gnd DFFSR_208/S FILL
XNAND2X1_1 BUFX2_12/Y AND2X2_2/Y DFFSR_28/gnd OAI22X1_7/D DFFSR_3/S NAND2X1
XFILL_0_NAND3X1_71 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_21_DFFSR_107 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_35_DFFSR_211 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_0_OAI21X1_117 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_0_AND2X2_21 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_11_DFFSR_110 OR2X2_3/gnd DFFSR_4/S FILL
XFILL_23_DFFPOSX1_47 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_25_DFFSR_214 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_1_XOR2X1_9 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_0_DFFSR_3 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_49_DFFSR_89 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_15_DFFSR_217 BUFX2_72/gnd DFFSR_201/S FILL
XINVX1_73 INVX1_73/A DFFSR_1/gnd INVX1_73/Y DFFSR_1/S INVX1
XFILL_5_DFFSR_86 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_7_DFFSR_104 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_22_DFFSR_79 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_33_DFFSR_39 INVX1_3/gnd DFFSR_79/S FILL
XFILL_48_DFFSR_135 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_8_NAND3X1_11 OR2X2_4/gnd DFFSR_32/S FILL
XINVX1_191 DFFSR_266/Q INVX1_67/gnd INVX1_191/Y DFFSR_175/S INVX1
XFILL_8_NAND3X1_184 BUFX2_8/gnd DFFSR_51/S FILL
XFILL_38_DFFSR_138 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_1_DFFSR_214 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_7_NAND3X1_14 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_18_3 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_4_BUFX2_24 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_28_DFFSR_141 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_1_NAND2X1_165 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_4_INVX1_188 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_33_2_0 INVX1_1/gnd DFFSR_53/S FILL
XFILL_42_DFFSR_245 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_6_NAND3X1_17 BUFX2_99/A DFFSR_7/S FILL
XFILL_4_CLKBUF1_9 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_18_DFFSR_144 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_14_NOR3X1_3 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_32_DFFSR_248 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_24_DFFSR_7 BUFX2_79/A DFFSR_7/S FILL
XFILL_5_NAND3X1_20 BUFX2_99/A DFFSR_7/S FILL
XFILL_22_DFFSR_251 BUFX2_7/gnd DFFSR_151/S FILL
XNAND3X1_17 DFFSR_59/D BUFX2_16/Y BUFX2_11/Y BUFX2_99/A NAND3X1_17/Y DFFSR_7/S NAND3X1
XFILL_4_NAND3X1_23 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_31_4_1 XOR2X1_4/gnd DFFSR_97/S FILL
XFILL_30_DFFSR_86 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_2_INVX1_80 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_41_DFFSR_46 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_3_NOR2X1_23 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_13_DFFPOSX1_22 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_3_NAND3X1_26 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_12_DFFSR_254 DFFSR_34/gnd DFFSR_1/S FILL
XDFFSR_144 DFFSR_200/D CLKBUF1_14/Y BUFX2_64/Y DFFSR_62/S DFFSR_144/D DFFSR_46/gnd
+ DFFSR_62/S DFFSR
XFILL_2_NAND3X1_29 OR2X2_4/gnd DFFSR_32/S FILL
XFILL_3_OAI22X1_11 BUFX2_99/A DFFSR_92/S FILL
XFILL_29_6_2 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_14_DFFSR_36 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_4_DFFSR_141 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_2_OAI22X1_14 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_1_BUFX2_71 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_1_NAND3X1_32 BUFX2_79/A DFFSR_7/S FILL
XFILL_45_DFFSR_172 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_8_DFFSR_248 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_0_NAND3X1_35 DFFSR_8/gnd DFFSR_8/S FILL
XFILL_1_OAI22X1_17 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_35_DFFSR_175 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_23_DFFPOSX1_11 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_49_DFFSR_279 BUFX2_99/A DFFSR_7/S FILL
XFILL_0_OAI22X1_20 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_45_DFFSR_3 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_25_DFFSR_178 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_49_DFFSR_53 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_38_DFFSR_93 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_15_DFFSR_181 INVX1_3/gnd DFFSR_79/S FILL
XFILL_7_NAND3X1_214 DFFSR_46/gnd DFFSR_62/S FILL
XFILL_3_DFFPOSX1_33 XOR2X1_4/gnd DFFSR_91/S FILL
XINVX1_37 INVX1_37/A BUFX2_77/gnd INVX1_37/Y DFFSR_98/S INVX1
XFILL_5_DFFSR_50 BUFX2_77/gnd DFFSR_5/S FILL
XDFFSR_90 DFFSR_98/D DFFSR_82/CLK DFFSR_35/R DFFSR_5/S DFFSR_82/Q BUFX2_77/gnd DFFSR_5/S
+ DFFSR
XFILL_22_DFFSR_43 BUFX2_98/A DFFSR_6/S FILL
XFILL_11_DFFSR_83 INVX1_3/gnd DFFSR_79/S FILL
XFILL_0_NOR2X1_60 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_2_OAI21X1_8 BUFX2_99/A DFFSR_7/S FILL
XINVX1_155 INVX1_155/A OR2X2_2/gnd INVX1_155/Y DFFSR_175/S INVX1
XFILL_38_DFFSR_102 DFFSR_4/gnd DFFSR_98/S FILL
XFILL_8_NAND3X1_148 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_1_DFFSR_178 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_0_INVX1_5 BUFX2_8/gnd DFFSR_81/S FILL
XFILL_1_7 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_28_DFFSR_105 INVX1_1/gnd DFFSR_53/S FILL
XFILL_1_NAND2X1_129 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_42_DFFSR_209 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_4_INVX1_152 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_7_AND2X2_19 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_18_DFFSR_108 OR2X2_6/gnd DFFSR_92/S FILL
XFILL_32_DFFSR_212 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_7_AND2X2_9 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_22_DFFSR_215 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_41_DFFSR_10 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_30_DFFSR_50 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_2_INVX1_44 OR2X2_4/gnd DFFSR_3/S FILL
XFILL_2_DFFSR_97 INVX1_1/gnd DFFSR_97/S FILL
XFILL_19_DFFSR_90 BUFX2_77/gnd DFFSR_5/S FILL
XFILL_39_1_2 BUFX2_79/A DFFSR_6/S FILL
XFILL_12_DFFSR_218 BUFX2_98/A DFFSR_32/S FILL
XFILL_22_DFFPOSX1_41 DFFSR_8/gnd DFFSR_60/S FILL
XDFFSR_108 DFFSR_116/D DFFSR_79/CLK DFFSR_7/R DFFSR_92/S DFFSR_100/Q OR2X2_6/gnd DFFSR_92/S
+ DFFSR
XFILL_4_DFFSR_105 INVX1_1/gnd DFFSR_53/S FILL
XFILL_6_NAND3X1_244 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_1_BUFX2_35 OR2X2_1/gnd DFFSR_59/S FILL
XFILL_45_DFFSR_136 NOR3X1_6/gnd DFFSR_79/S FILL
XFILL_8_DFFSR_212 OR2X2_2/gnd DFFSR_175/S FILL
XFILL_35_DFFSR_139 DFFSR_34/gnd DFFSR_34/S FILL
XFILL_49_DFFSR_243 BUFX2_7/gnd DFFSR_151/S FILL
XFILL_9_OAI21X1_100 INVX1_3/gnd DFFSR_79/S FILL
XFILL_11_DFFSR_1 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_25_DFFSR_142 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_49_DFFSR_17 DFFSR_28/gnd DFFSR_3/S FILL
XFILL_1_INVX1_189 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_39_DFFSR_246 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_38_DFFSR_57 BUFX2_79/A DFFSR_6/S FILL
XFILL_27_DFFSR_97 INVX1_1/gnd DFFSR_97/S FILL
XFILL_15_DFFSR_145 BUFX2_72/gnd DFFSR_201/S FILL
XFILL_7_NAND3X1_178 NOR3X1_6/gnd DFFSR_91/S FILL
XFILL_29_DFFSR_249 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_0_NAND2X1_159 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_19_DFFSR_252 AND2X2_38/B DFFSR_23/S FILL
XDFFSR_54 DFFSR_54/Q AOI21X1_3/B DFFSR_1/R DFFSR_54/S DFFSR_62/Q INVX1_39/gnd DFFSR_54/S
+ DFFSR
XFILL_5_DFFSR_14 INVX1_1/gnd DFFSR_53/S FILL
XFILL_11_DFFSR_47 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_0_NOR2X1_24 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_8_NAND3X1_112 DFFSR_1/gnd DFFSR_1/S FILL
XINVX1_119 BUFX2_39/Y DFFSR_46/gnd INVX1_119/Y DFFSR_54/S INVX1
XFILL_1_DFFSR_142 XOR2X1_1/gnd DFFSR_151/S FILL
XFILL_12_DFFPOSX1_16 INVX1_67/gnd DFFSR_175/S FILL
XFILL_4_INVX1_116 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_42_DFFSR_173 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_46_DFFSR_64 OR2X2_3/gnd DFFSR_60/S FILL
XFILL_5_DFFSR_249 BUFX2_72/gnd DFFSR_276/S FILL
XFILL_32_DFFSR_176 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_46_DFFSR_280 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_22_DFFSR_179 OR2X2_1/gnd DFFSR_51/S FILL
XFILL_2_DFFSR_61 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_30_DFFSR_14 INVX1_1/gnd DFFSR_53/S FILL
XFILL_19_DFFSR_54 INVX1_39/gnd DFFSR_54/S FILL
XFILL_12_DFFSR_182 XOR2X1_1/gnd DFFSR_208/S FILL
XFILL_6_BUFX2_89 INVX1_1/gnd DFFSR_97/S FILL
XFILL_20_CLKBUF1_44 DFFSR_1/gnd DFFSR_81/S FILL
XFILL_6_NAND3X1_208 DFFSR_46/gnd DFFSR_54/S FILL
XFILL_45_DFFSR_100 INVX1_1/gnd DFFSR_97/S FILL
XFILL_19_CLKBUF1_47 BUFX2_98/A DFFSR_32/S FILL
XFILL_8_DFFSR_176 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_2_DFFPOSX1_27 DFFSR_34/gnd DFFSR_1/S FILL
XFILL_35_DFFSR_103 DFFSR_8/gnd DFFSR_60/S FILL
XAND2X2_23 AND2X2_23/A AND2X2_23/B OR2X2_1/gnd AND2X2_23/Y DFFSR_59/S AND2X2
XFILL_49_DFFSR_207 DFFSR_62/gnd DFFSR_62/S FILL
XNAND3X1_244 INVX1_170/Y AOI21X1_45/B AOI21X1_45/A DFFSR_28/gnd NAND2X1_113/B DFFSR_8/S
+ NAND3X1
XFILL_25_DFFSR_106 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_1_INVX1_153 INVX1_67/gnd DFFSR_175/S FILL
XFILL_39_DFFSR_210 BUFX2_98/A DFFSR_6/S FILL
XFILL_27_DFFSR_61 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_38_DFFSR_21 DFFSR_5/gnd DFFSR_5/S FILL
XFILL_4_AND2X2_20 OR2X2_6/gnd DFFSR_53/S FILL
XFILL_15_DFFSR_109 DFFSR_4/gnd DFFSR_4/S FILL
XFILL_7_NAND3X1_142 INVX1_67/gnd DFFSR_175/S FILL
XFILL_29_DFFSR_213 INVX1_3/gnd DFFSR_23/S FILL
XFILL_11_DFFPOSX1_46 INVX1_39/gnd DFFSR_34/S FILL
XFILL_19_DFFSR_216 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_0_NAND2X1_123 BUFX2_77/gnd DFFSR_98/S FILL
XDFFSR_18 DFFSR_34/D DFFSR_79/CLK DFFSR_7/R DFFSR_91/S DFFSR_18/D NOR3X1_6/gnd DFFSR_91/S
+ DFFSR
XFILL_11_DFFSR_11 DFFSR_1/gnd DFFSR_1/S FILL
XFILL_1_DFFSR_106 XOR2X1_4/gnd DFFSR_91/S FILL
XFILL_21_DFFPOSX1_35 INVX1_39/gnd DFFSR_54/S FILL
XFILL_42_DFFSR_137 BUFX2_7/gnd DFFSR_216/S FILL
XFILL_46_DFFSR_28 DFFSR_28/gnd DFFSR_8/S FILL
XFILL_35_DFFSR_68 BUFX2_98/A DFFSR_6/S FILL
XFILL_5_DFFSR_213 INVX1_3/gnd DFFSR_23/S FILL
XFILL_32_DFFSR_140 DFFSR_62/gnd DFFSR_208/S FILL
XFILL_5_NAND3X1_238 BUFX2_77/gnd DFFSR_98/S FILL
XFILL_46_DFFSR_244 DFFSR_1/gnd DFFSR_81/S FILL
.ends


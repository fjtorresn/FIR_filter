module fir2n (clk, rst, din, dout);

input clk;
input rst;
input [7:0] din;
output [7:0] dout;

wire vdd = 1'b1;
wire gnd = 1'b0;

BUFX2 BUFX2_1 ( .A(clk2_clkout), .Y(clk2_clkout_hier0_bF_buf5) );
BUFX2 BUFX2_2 ( .A(clk2_clkout), .Y(clk2_clkout_hier0_bF_buf4) );
BUFX2 BUFX2_3 ( .A(clk2_clkout), .Y(clk2_clkout_hier0_bF_buf3) );
BUFX2 BUFX2_4 ( .A(clk2_clkout), .Y(clk2_clkout_hier0_bF_buf2) );
BUFX2 BUFX2_5 ( .A(clk2_clkout), .Y(clk2_clkout_hier0_bF_buf1) );
BUFX2 BUFX2_6 ( .A(clk2_clkout), .Y(clk2_clkout_hier0_bF_buf0) );
BUFX2 BUFX2_7 ( .A(counterup_counter_0_), .Y(counterup_counter_0_bF_buf3_) );
BUFX2 BUFX2_8 ( .A(counterup_counter_0_), .Y(counterup_counter_0_bF_buf2_) );
BUFX2 BUFX2_9 ( .A(counterup_counter_0_), .Y(counterup_counter_0_bF_buf1_) );
BUFX2 BUFX2_10 ( .A(counterup_counter_0_), .Y(counterup_counter_0_bF_buf0_) );
CLKBUF1 CLKBUF1_1 ( .A(clk2_clkout_hier0_bF_buf5), .Y(clk2_clkout_bF_buf41) );
CLKBUF1 CLKBUF1_2 ( .A(clk2_clkout_hier0_bF_buf4), .Y(clk2_clkout_bF_buf40) );
CLKBUF1 CLKBUF1_3 ( .A(clk2_clkout_hier0_bF_buf3), .Y(clk2_clkout_bF_buf39) );
CLKBUF1 CLKBUF1_4 ( .A(clk2_clkout_hier0_bF_buf2), .Y(clk2_clkout_bF_buf38) );
CLKBUF1 CLKBUF1_5 ( .A(clk2_clkout_hier0_bF_buf1), .Y(clk2_clkout_bF_buf37) );
CLKBUF1 CLKBUF1_6 ( .A(clk2_clkout_hier0_bF_buf0), .Y(clk2_clkout_bF_buf36) );
CLKBUF1 CLKBUF1_7 ( .A(clk2_clkout_hier0_bF_buf5), .Y(clk2_clkout_bF_buf35) );
CLKBUF1 CLKBUF1_8 ( .A(clk2_clkout_hier0_bF_buf4), .Y(clk2_clkout_bF_buf34) );
CLKBUF1 CLKBUF1_9 ( .A(clk2_clkout_hier0_bF_buf3), .Y(clk2_clkout_bF_buf33) );
CLKBUF1 CLKBUF1_10 ( .A(clk2_clkout_hier0_bF_buf2), .Y(clk2_clkout_bF_buf32) );
CLKBUF1 CLKBUF1_11 ( .A(clk2_clkout_hier0_bF_buf1), .Y(clk2_clkout_bF_buf31) );
CLKBUF1 CLKBUF1_12 ( .A(clk2_clkout_hier0_bF_buf0), .Y(clk2_clkout_bF_buf30) );
CLKBUF1 CLKBUF1_13 ( .A(clk2_clkout_hier0_bF_buf5), .Y(clk2_clkout_bF_buf29) );
CLKBUF1 CLKBUF1_14 ( .A(clk2_clkout_hier0_bF_buf4), .Y(clk2_clkout_bF_buf28) );
CLKBUF1 CLKBUF1_15 ( .A(clk2_clkout_hier0_bF_buf3), .Y(clk2_clkout_bF_buf27) );
CLKBUF1 CLKBUF1_16 ( .A(clk2_clkout_hier0_bF_buf2), .Y(clk2_clkout_bF_buf26) );
CLKBUF1 CLKBUF1_17 ( .A(clk2_clkout_hier0_bF_buf1), .Y(clk2_clkout_bF_buf25) );
CLKBUF1 CLKBUF1_18 ( .A(clk2_clkout_hier0_bF_buf0), .Y(clk2_clkout_bF_buf24) );
CLKBUF1 CLKBUF1_19 ( .A(clk2_clkout_hier0_bF_buf5), .Y(clk2_clkout_bF_buf23) );
CLKBUF1 CLKBUF1_20 ( .A(clk2_clkout_hier0_bF_buf4), .Y(clk2_clkout_bF_buf22) );
CLKBUF1 CLKBUF1_21 ( .A(clk2_clkout_hier0_bF_buf3), .Y(clk2_clkout_bF_buf21) );
CLKBUF1 CLKBUF1_22 ( .A(clk2_clkout_hier0_bF_buf2), .Y(clk2_clkout_bF_buf20) );
CLKBUF1 CLKBUF1_23 ( .A(clk2_clkout_hier0_bF_buf1), .Y(clk2_clkout_bF_buf19) );
CLKBUF1 CLKBUF1_24 ( .A(clk2_clkout_hier0_bF_buf0), .Y(clk2_clkout_bF_buf18) );
CLKBUF1 CLKBUF1_25 ( .A(clk2_clkout_hier0_bF_buf5), .Y(clk2_clkout_bF_buf17) );
CLKBUF1 CLKBUF1_26 ( .A(clk2_clkout_hier0_bF_buf4), .Y(clk2_clkout_bF_buf16) );
CLKBUF1 CLKBUF1_27 ( .A(clk2_clkout_hier0_bF_buf3), .Y(clk2_clkout_bF_buf15) );
CLKBUF1 CLKBUF1_28 ( .A(clk2_clkout_hier0_bF_buf2), .Y(clk2_clkout_bF_buf14) );
CLKBUF1 CLKBUF1_29 ( .A(clk2_clkout_hier0_bF_buf1), .Y(clk2_clkout_bF_buf13) );
CLKBUF1 CLKBUF1_30 ( .A(clk2_clkout_hier0_bF_buf0), .Y(clk2_clkout_bF_buf12) );
CLKBUF1 CLKBUF1_31 ( .A(clk2_clkout_hier0_bF_buf5), .Y(clk2_clkout_bF_buf11) );
CLKBUF1 CLKBUF1_32 ( .A(clk2_clkout_hier0_bF_buf4), .Y(clk2_clkout_bF_buf10) );
CLKBUF1 CLKBUF1_33 ( .A(clk2_clkout_hier0_bF_buf3), .Y(clk2_clkout_bF_buf9) );
CLKBUF1 CLKBUF1_34 ( .A(clk2_clkout_hier0_bF_buf2), .Y(clk2_clkout_bF_buf8) );
CLKBUF1 CLKBUF1_35 ( .A(clk2_clkout_hier0_bF_buf1), .Y(clk2_clkout_bF_buf7) );
CLKBUF1 CLKBUF1_36 ( .A(clk2_clkout_hier0_bF_buf0), .Y(clk2_clkout_bF_buf6) );
CLKBUF1 CLKBUF1_37 ( .A(clk2_clkout_hier0_bF_buf5), .Y(clk2_clkout_bF_buf5) );
CLKBUF1 CLKBUF1_38 ( .A(clk2_clkout_hier0_bF_buf4), .Y(clk2_clkout_bF_buf4) );
CLKBUF1 CLKBUF1_39 ( .A(clk2_clkout_hier0_bF_buf3), .Y(clk2_clkout_bF_buf3) );
CLKBUF1 CLKBUF1_40 ( .A(clk2_clkout_hier0_bF_buf2), .Y(clk2_clkout_bF_buf2) );
CLKBUF1 CLKBUF1_41 ( .A(clk2_clkout_hier0_bF_buf1), .Y(clk2_clkout_bF_buf1) );
CLKBUF1 CLKBUF1_42 ( .A(clk2_clkout_hier0_bF_buf0), .Y(clk2_clkout_bF_buf0) );
BUFX2 BUFX2_11 ( .A(_4_), .Y(_4__bF_buf3) );
BUFX2 BUFX2_12 ( .A(_4_), .Y(_4__bF_buf2) );
BUFX2 BUFX2_13 ( .A(_4_), .Y(_4__bF_buf1) );
BUFX2 BUFX2_14 ( .A(_4_), .Y(_4__bF_buf0) );
CLKBUF1 CLKBUF1_43 ( .A(clk), .Y(clk_bF_buf6) );
CLKBUF1 CLKBUF1_44 ( .A(clk), .Y(clk_bF_buf5) );
CLKBUF1 CLKBUF1_45 ( .A(clk), .Y(clk_bF_buf4) );
CLKBUF1 CLKBUF1_46 ( .A(clk), .Y(clk_bF_buf3) );
CLKBUF1 CLKBUF1_47 ( .A(clk), .Y(clk_bF_buf2) );
CLKBUF1 CLKBUF1_48 ( .A(clk), .Y(clk_bF_buf1) );
CLKBUF1 CLKBUF1_49 ( .A(clk), .Y(clk_bF_buf0) );
BUFX2 BUFX2_15 ( .A(_36_), .Y(_36__bF_buf3) );
BUFX2 BUFX2_16 ( .A(_36_), .Y(_36__bF_buf2) );
BUFX2 BUFX2_17 ( .A(_36_), .Y(_36__bF_buf1) );
BUFX2 BUFX2_18 ( .A(_36_), .Y(_36__bF_buf0) );
BUFX2 BUFX2_19 ( .A(_33_), .Y(_33__bF_buf3) );
BUFX2 BUFX2_20 ( .A(_33_), .Y(_33__bF_buf2) );
BUFX2 BUFX2_21 ( .A(_33_), .Y(_33__bF_buf1) );
BUFX2 BUFX2_22 ( .A(_33_), .Y(_33__bF_buf0) );
BUFX2 BUFX2_23 ( .A(_229_), .Y(_229__bF_buf3) );
BUFX2 BUFX2_24 ( .A(_229_), .Y(_229__bF_buf2) );
BUFX2 BUFX2_25 ( .A(_229_), .Y(_229__bF_buf1) );
BUFX2 BUFX2_26 ( .A(_229_), .Y(_229__bF_buf0) );
BUFX2 BUFX2_27 ( .A(_261_), .Y(_261__bF_buf3) );
BUFX2 BUFX2_28 ( .A(_261_), .Y(_261__bF_buf2) );
BUFX2 BUFX2_29 ( .A(_261_), .Y(_261__bF_buf1) );
BUFX2 BUFX2_30 ( .A(_261_), .Y(_261__bF_buf0) );
BUFX2 BUFX2_31 ( .A(_258_), .Y(_258__bF_buf3) );
BUFX2 BUFX2_32 ( .A(_258_), .Y(_258__bF_buf2) );
BUFX2 BUFX2_33 ( .A(_258_), .Y(_258__bF_buf1) );
BUFX2 BUFX2_34 ( .A(_258_), .Y(_258__bF_buf0) );
BUFX2 BUFX2_35 ( .A(rst), .Y(rst_bF_buf5) );
BUFX2 BUFX2_36 ( .A(rst), .Y(rst_bF_buf4) );
BUFX2 BUFX2_37 ( .A(rst), .Y(rst_bF_buf3) );
BUFX2 BUFX2_38 ( .A(rst), .Y(rst_bF_buf2) );
BUFX2 BUFX2_39 ( .A(rst), .Y(rst_bF_buf1) );
BUFX2 BUFX2_40 ( .A(rst), .Y(rst_bF_buf0) );
BUFX2 BUFX2_41 ( .A(_0_), .Y(_0__bF_buf10) );
BUFX2 BUFX2_42 ( .A(_0_), .Y(_0__bF_buf9) );
BUFX2 BUFX2_43 ( .A(_0_), .Y(_0__bF_buf8) );
BUFX2 BUFX2_44 ( .A(_0_), .Y(_0__bF_buf7) );
BUFX2 BUFX2_45 ( .A(_0_), .Y(_0__bF_buf6) );
BUFX2 BUFX2_46 ( .A(_0_), .Y(_0__bF_buf5) );
BUFX2 BUFX2_47 ( .A(_0_), .Y(_0__bF_buf4) );
BUFX2 BUFX2_48 ( .A(_0_), .Y(_0__bF_buf3) );
BUFX2 BUFX2_49 ( .A(_0_), .Y(_0__bF_buf2) );
BUFX2 BUFX2_50 ( .A(_0_), .Y(_0__bF_buf1) );
BUFX2 BUFX2_51 ( .A(_0_), .Y(_0__bF_buf0) );
BUFX2 BUFX2_52 ( .A(mac1_reset), .Y(mac1_reset_bF_buf3) );
BUFX2 BUFX2_53 ( .A(mac1_reset), .Y(mac1_reset_bF_buf2) );
BUFX2 BUFX2_54 ( .A(mac1_reset), .Y(mac1_reset_bF_buf1) );
BUFX2 BUFX2_55 ( .A(mac1_reset), .Y(mac1_reset_bF_buf0) );
BUFX2 BUFX2_56 ( .A(rom1_data_0_), .Y(rom1_data_0_bF_buf3_) );
BUFX2 BUFX2_57 ( .A(rom1_data_0_), .Y(rom1_data_0_bF_buf2_) );
BUFX2 BUFX2_58 ( .A(rom1_data_0_), .Y(rom1_data_0_bF_buf1_) );
BUFX2 BUFX2_59 ( .A(rom1_data_0_), .Y(rom1_data_0_bF_buf0_) );
BUFX2 BUFX2_60 ( .A(_225_), .Y(_225__bF_buf10) );
BUFX2 BUFX2_61 ( .A(_225_), .Y(_225__bF_buf9) );
BUFX2 BUFX2_62 ( .A(_225_), .Y(_225__bF_buf8) );
BUFX2 BUFX2_63 ( .A(_225_), .Y(_225__bF_buf7) );
BUFX2 BUFX2_64 ( .A(_225_), .Y(_225__bF_buf6) );
BUFX2 BUFX2_65 ( .A(_225_), .Y(_225__bF_buf5) );
BUFX2 BUFX2_66 ( .A(_225_), .Y(_225__bF_buf4) );
BUFX2 BUFX2_67 ( .A(_225_), .Y(_225__bF_buf3) );
BUFX2 BUFX2_68 ( .A(_225_), .Y(_225__bF_buf2) );
BUFX2 BUFX2_69 ( .A(_225_), .Y(_225__bF_buf1) );
BUFX2 BUFX2_70 ( .A(_225_), .Y(_225__bF_buf0) );
BUFX2 BUFX2_71 ( .A(reg3_dataout_0_), .Y(dout[0]) );
BUFX2 BUFX2_72 ( .A(reg3_dataout_1_), .Y(dout[1]) );
BUFX2 BUFX2_73 ( .A(reg3_dataout_2_), .Y(dout[2]) );
BUFX2 BUFX2_74 ( .A(reg3_dataout_3_), .Y(dout[3]) );
BUFX2 BUFX2_75 ( .A(reg3_dataout_4_), .Y(dout[4]) );
BUFX2 BUFX2_76 ( .A(reg3_dataout_5_), .Y(dout[5]) );
BUFX2 BUFX2_77 ( .A(reg3_dataout_6_), .Y(dout[6]) );
BUFX2 BUFX2_78 ( .A(reg3_dataout_7_), .Y(dout[7]) );
INVX1 INVX1_1 ( .A(asr1_rom_6__0_), .Y(_1_) );
INVX1 INVX1_2 ( .A(asr1_rom_5__0_), .Y(_2_) );
INVX1 INVX1_3 ( .A(counterup_counter_3_), .Y(_3_) );
AND2X2 AND2X2_1 ( .A(_3_), .B(counterup_counter_2_), .Y(_4_) );
INVX1 INVX1_4 ( .A(counterup_counter_1_), .Y(_5_) );
AND2X2 AND2X2_2 ( .A(_5_), .B(counterup_counter_0_bF_buf3_), .Y(_6_) );
NAND2X1 NAND2X1_1 ( .A(_4__bF_buf3), .B(_6_), .Y(_7_) );
NOR2X1 NOR2X1_1 ( .A(counterup_counter_0_bF_buf2_), .B(_5_), .Y(_8_) );
NAND2X1 NAND2X1_2 ( .A(_8_), .B(_4__bF_buf2), .Y(_9_) );
OAI22X1 OAI22X1_1 ( .A(_1_), .B(_9_), .C(_2_), .D(_7_), .Y(_10_) );
INVX1 INVX1_5 ( .A(asr1_rom_10__0_), .Y(_11_) );
INVX1 INVX1_6 ( .A(asr1_rom_9__0_), .Y(_12_) );
NOR2X1 NOR2X1_2 ( .A(counterup_counter_2_), .B(_3_), .Y(_13_) );
NAND2X1 NAND2X1_3 ( .A(_13_), .B(_6_), .Y(_14_) );
NAND2X1 NAND2X1_4 ( .A(_8_), .B(_13_), .Y(_15_) );
OAI22X1 OAI22X1_2 ( .A(_11_), .B(_15_), .C(_12_), .D(_14_), .Y(_16_) );
NOR2X1 NOR2X1_3 ( .A(_16_), .B(_10_), .Y(_17_) );
INVX1 INVX1_7 ( .A(asr1_rom_2__0_), .Y(_18_) );
INVX1 INVX1_8 ( .A(asr1_rom_1__0_), .Y(_19_) );
NOR2X1 NOR2X1_4 ( .A(counterup_counter_3_), .B(counterup_counter_2_), .Y(_20_) );
NAND2X1 NAND2X1_5 ( .A(_20_), .B(_6_), .Y(_21_) );
NAND2X1 NAND2X1_6 ( .A(_20_), .B(_8_), .Y(_22_) );
OAI22X1 OAI22X1_3 ( .A(_18_), .B(_22_), .C(_19_), .D(_21_), .Y(_23_) );
INVX1 INVX1_9 ( .A(asr1_rom_14__0_), .Y(_24_) );
NAND2X1 NAND2X1_7 ( .A(counterup_counter_0_bF_buf1_), .B(_5_), .Y(_25_) );
NAND2X1 NAND2X1_8 ( .A(counterup_counter_3_), .B(counterup_counter_2_), .Y(_26_) );
NOR2X1 NOR2X1_5 ( .A(_26_), .B(_25_), .Y(_27_) );
NAND2X1 NAND2X1_9 ( .A(asr1_rom_13__0_), .B(_27_), .Y(_28_) );
AND2X2 AND2X2_3 ( .A(counterup_counter_3_), .B(counterup_counter_2_), .Y(_29_) );
NAND2X1 NAND2X1_10 ( .A(_29_), .B(_8_), .Y(_30_) );
OAI21X1 OAI21X1_1 ( .A(_24_), .B(_30_), .C(_28_), .Y(_31_) );
NOR2X1 NOR2X1_6 ( .A(_23_), .B(_31_), .Y(_32_) );
AND2X2 AND2X2_4 ( .A(counterup_counter_1_), .B(counterup_counter_0_bF_buf0_), .Y(_33_) );
AND2X2 AND2X2_5 ( .A(_33__bF_buf3), .B(_20_), .Y(_34_) );
NAND2X1 NAND2X1_11 ( .A(asr1_rom_3__0_), .B(_34_), .Y(_35_) );
NOR2X1 NOR2X1_7 ( .A(counterup_counter_1_), .B(counterup_counter_0_bF_buf3_), .Y(_36_) );
NAND3X1 NAND3X1_1 ( .A(asr1_rom_4__0_), .B(_36__bF_buf3), .C(_4__bF_buf1), .Y(_37_) );
NAND3X1 NAND3X1_2 ( .A(asr1_rom_0__0_), .B(_20_), .C(_36__bF_buf2), .Y(_38_) );
NAND3X1 NAND3X1_3 ( .A(asr1_en_0_), .B(_29_), .C(_33__bF_buf2), .Y(_39_) );
AND2X2 AND2X2_6 ( .A(_39_), .B(_38_), .Y(_40_) );
NAND3X1 NAND3X1_4 ( .A(_35_), .B(_37_), .C(_40_), .Y(_41_) );
NAND3X1 NAND3X1_5 ( .A(asr1_rom_7__0_), .B(_33__bF_buf1), .C(_4__bF_buf0), .Y(_42_) );
NAND3X1 NAND3X1_6 ( .A(asr1_rom_8__0_), .B(_36__bF_buf1), .C(_13_), .Y(_43_) );
NAND2X1 NAND2X1_12 ( .A(counterup_counter_1_), .B(counterup_counter_0_bF_buf2_), .Y(_44_) );
NOR3X1 NOR3X1_1 ( .A(counterup_counter_2_), .B(_3_), .C(_44_), .Y(_45_) );
NOR3X1 NOR3X1_2 ( .A(counterup_counter_1_), .B(counterup_counter_0_bF_buf1_), .C(_26_), .Y(_46_) );
AOI22X1 AOI22X1_1 ( .A(_46_), .B(asr1_rom_12__0_), .C(asr1_rom_11__0_), .D(_45_), .Y(_47_) );
NAND3X1 NAND3X1_7 ( .A(_42_), .B(_43_), .C(_47_), .Y(_48_) );
NOR2X1 NOR2X1_8 ( .A(_41_), .B(_48_), .Y(_49_) );
NAND3X1 NAND3X1_8 ( .A(_17_), .B(_32_), .C(_49_), .Y(asr1_dataout_0_) );
INVX1 INVX1_10 ( .A(asr1_rom_6__1_), .Y(_50_) );
INVX1 INVX1_11 ( .A(asr1_rom_5__1_), .Y(_51_) );
OAI22X1 OAI22X1_4 ( .A(_50_), .B(_9_), .C(_51_), .D(_7_), .Y(_52_) );
INVX1 INVX1_12 ( .A(asr1_rom_10__1_), .Y(_53_) );
INVX1 INVX1_13 ( .A(asr1_rom_9__1_), .Y(_54_) );
OAI22X1 OAI22X1_5 ( .A(_53_), .B(_15_), .C(_54_), .D(_14_), .Y(_55_) );
NOR2X1 NOR2X1_9 ( .A(_55_), .B(_52_), .Y(_56_) );
INVX1 INVX1_14 ( .A(asr1_rom_2__1_), .Y(_57_) );
INVX1 INVX1_15 ( .A(asr1_rom_1__1_), .Y(_58_) );
OAI22X1 OAI22X1_6 ( .A(_57_), .B(_22_), .C(_58_), .D(_21_), .Y(_59_) );
INVX1 INVX1_16 ( .A(asr1_rom_14__1_), .Y(_60_) );
NAND2X1 NAND2X1_13 ( .A(asr1_rom_13__1_), .B(_27_), .Y(_61_) );
OAI21X1 OAI21X1_2 ( .A(_60_), .B(_30_), .C(_61_), .Y(_62_) );
NOR2X1 NOR2X1_10 ( .A(_59_), .B(_62_), .Y(_63_) );
NAND2X1 NAND2X1_14 ( .A(asr1_rom_3__1_), .B(_34_), .Y(_64_) );
NAND3X1 NAND3X1_9 ( .A(asr1_rom_4__1_), .B(_36__bF_buf0), .C(_4__bF_buf3), .Y(_65_) );
NAND3X1 NAND3X1_10 ( .A(asr1_rom_0__1_), .B(_20_), .C(_36__bF_buf3), .Y(_66_) );
NAND3X1 NAND3X1_11 ( .A(asr1_en_1_), .B(_29_), .C(_33__bF_buf0), .Y(_67_) );
AND2X2 AND2X2_7 ( .A(_67_), .B(_66_), .Y(_68_) );
NAND3X1 NAND3X1_12 ( .A(_64_), .B(_65_), .C(_68_), .Y(_69_) );
NAND3X1 NAND3X1_13 ( .A(asr1_rom_7__1_), .B(_33__bF_buf3), .C(_4__bF_buf2), .Y(_70_) );
NAND3X1 NAND3X1_14 ( .A(asr1_rom_8__1_), .B(_36__bF_buf2), .C(_13_), .Y(_71_) );
AOI22X1 AOI22X1_2 ( .A(_46_), .B(asr1_rom_12__1_), .C(asr1_rom_11__1_), .D(_45_), .Y(_72_) );
NAND3X1 NAND3X1_15 ( .A(_70_), .B(_71_), .C(_72_), .Y(_73_) );
NOR2X1 NOR2X1_11 ( .A(_69_), .B(_73_), .Y(_74_) );
NAND3X1 NAND3X1_16 ( .A(_56_), .B(_63_), .C(_74_), .Y(asr1_dataout_1_) );
INVX1 INVX1_17 ( .A(asr1_rom_6__2_), .Y(_75_) );
INVX1 INVX1_18 ( .A(asr1_rom_5__2_), .Y(_76_) );
OAI22X1 OAI22X1_7 ( .A(_75_), .B(_9_), .C(_76_), .D(_7_), .Y(_77_) );
INVX1 INVX1_19 ( .A(asr1_rom_10__2_), .Y(_78_) );
INVX1 INVX1_20 ( .A(asr1_rom_9__2_), .Y(_79_) );
OAI22X1 OAI22X1_8 ( .A(_78_), .B(_15_), .C(_79_), .D(_14_), .Y(_80_) );
NOR2X1 NOR2X1_12 ( .A(_80_), .B(_77_), .Y(_81_) );
INVX1 INVX1_21 ( .A(asr1_rom_2__2_), .Y(_82_) );
INVX1 INVX1_22 ( .A(asr1_rom_1__2_), .Y(_83_) );
OAI22X1 OAI22X1_9 ( .A(_82_), .B(_22_), .C(_83_), .D(_21_), .Y(_84_) );
INVX1 INVX1_23 ( .A(asr1_rom_14__2_), .Y(_85_) );
NAND2X1 NAND2X1_15 ( .A(asr1_rom_13__2_), .B(_27_), .Y(_86_) );
OAI21X1 OAI21X1_3 ( .A(_85_), .B(_30_), .C(_86_), .Y(_87_) );
NOR2X1 NOR2X1_13 ( .A(_84_), .B(_87_), .Y(_88_) );
NAND2X1 NAND2X1_16 ( .A(asr1_rom_3__2_), .B(_34_), .Y(_89_) );
NAND3X1 NAND3X1_17 ( .A(asr1_rom_4__2_), .B(_36__bF_buf1), .C(_4__bF_buf1), .Y(_90_) );
NAND3X1 NAND3X1_18 ( .A(asr1_rom_0__2_), .B(_20_), .C(_36__bF_buf0), .Y(_91_) );
NAND3X1 NAND3X1_19 ( .A(asr1_en_2_), .B(_29_), .C(_33__bF_buf2), .Y(_92_) );
AND2X2 AND2X2_8 ( .A(_92_), .B(_91_), .Y(_93_) );
NAND3X1 NAND3X1_20 ( .A(_89_), .B(_90_), .C(_93_), .Y(_94_) );
NAND3X1 NAND3X1_21 ( .A(asr1_rom_7__2_), .B(_33__bF_buf1), .C(_4__bF_buf0), .Y(_95_) );
NAND3X1 NAND3X1_22 ( .A(asr1_rom_8__2_), .B(_36__bF_buf3), .C(_13_), .Y(_96_) );
AOI22X1 AOI22X1_3 ( .A(_46_), .B(asr1_rom_12__2_), .C(asr1_rom_11__2_), .D(_45_), .Y(_97_) );
NAND3X1 NAND3X1_23 ( .A(_95_), .B(_96_), .C(_97_), .Y(_98_) );
NOR2X1 NOR2X1_14 ( .A(_94_), .B(_98_), .Y(_99_) );
NAND3X1 NAND3X1_24 ( .A(_81_), .B(_88_), .C(_99_), .Y(asr1_dataout_2_) );
INVX1 INVX1_24 ( .A(asr1_rom_6__3_), .Y(_100_) );
INVX1 INVX1_25 ( .A(asr1_rom_5__3_), .Y(_101_) );
OAI22X1 OAI22X1_10 ( .A(_100_), .B(_9_), .C(_101_), .D(_7_), .Y(_102_) );
INVX1 INVX1_26 ( .A(asr1_rom_10__3_), .Y(_103_) );
INVX1 INVX1_27 ( .A(asr1_rom_9__3_), .Y(_104_) );
OAI22X1 OAI22X1_11 ( .A(_103_), .B(_15_), .C(_104_), .D(_14_), .Y(_105_) );
NOR2X1 NOR2X1_15 ( .A(_105_), .B(_102_), .Y(_106_) );
INVX1 INVX1_28 ( .A(asr1_rom_2__3_), .Y(_107_) );
INVX1 INVX1_29 ( .A(asr1_rom_1__3_), .Y(_108_) );
OAI22X1 OAI22X1_12 ( .A(_107_), .B(_22_), .C(_108_), .D(_21_), .Y(_109_) );
INVX1 INVX1_30 ( .A(asr1_rom_14__3_), .Y(_110_) );
NAND2X1 NAND2X1_17 ( .A(asr1_rom_13__3_), .B(_27_), .Y(_111_) );
OAI21X1 OAI21X1_4 ( .A(_110_), .B(_30_), .C(_111_), .Y(_112_) );
NOR2X1 NOR2X1_16 ( .A(_109_), .B(_112_), .Y(_113_) );
NAND2X1 NAND2X1_18 ( .A(asr1_rom_3__3_), .B(_34_), .Y(_114_) );
NAND3X1 NAND3X1_25 ( .A(asr1_rom_4__3_), .B(_36__bF_buf2), .C(_4__bF_buf3), .Y(_115_) );
NAND3X1 NAND3X1_26 ( .A(asr1_rom_0__3_), .B(_20_), .C(_36__bF_buf1), .Y(_116_) );
NAND3X1 NAND3X1_27 ( .A(asr1_en_3_), .B(_29_), .C(_33__bF_buf0), .Y(_117_) );
AND2X2 AND2X2_9 ( .A(_117_), .B(_116_), .Y(_118_) );
NAND3X1 NAND3X1_28 ( .A(_114_), .B(_115_), .C(_118_), .Y(_119_) );
NAND3X1 NAND3X1_29 ( .A(asr1_rom_7__3_), .B(_33__bF_buf3), .C(_4__bF_buf2), .Y(_120_) );
NAND3X1 NAND3X1_30 ( .A(asr1_rom_8__3_), .B(_36__bF_buf0), .C(_13_), .Y(_121_) );
AOI22X1 AOI22X1_4 ( .A(_46_), .B(asr1_rom_12__3_), .C(asr1_rom_11__3_), .D(_45_), .Y(_122_) );
NAND3X1 NAND3X1_31 ( .A(_120_), .B(_121_), .C(_122_), .Y(_123_) );
NOR2X1 NOR2X1_17 ( .A(_119_), .B(_123_), .Y(_124_) );
NAND3X1 NAND3X1_32 ( .A(_106_), .B(_113_), .C(_124_), .Y(asr1_dataout_3_) );
INVX1 INVX1_31 ( .A(asr1_rom_6__4_), .Y(_125_) );
INVX1 INVX1_32 ( .A(asr1_rom_5__4_), .Y(_126_) );
OAI22X1 OAI22X1_13 ( .A(_125_), .B(_9_), .C(_126_), .D(_7_), .Y(_127_) );
INVX1 INVX1_33 ( .A(asr1_rom_10__4_), .Y(_128_) );
INVX1 INVX1_34 ( .A(asr1_rom_9__4_), .Y(_129_) );
OAI22X1 OAI22X1_14 ( .A(_128_), .B(_15_), .C(_129_), .D(_14_), .Y(_130_) );
NOR2X1 NOR2X1_18 ( .A(_130_), .B(_127_), .Y(_131_) );
INVX1 INVX1_35 ( .A(asr1_rom_2__4_), .Y(_132_) );
INVX1 INVX1_36 ( .A(asr1_rom_1__4_), .Y(_133_) );
OAI22X1 OAI22X1_15 ( .A(_132_), .B(_22_), .C(_133_), .D(_21_), .Y(_134_) );
INVX1 INVX1_37 ( .A(asr1_rom_14__4_), .Y(_135_) );
NAND2X1 NAND2X1_19 ( .A(asr1_rom_13__4_), .B(_27_), .Y(_136_) );
OAI21X1 OAI21X1_5 ( .A(_135_), .B(_30_), .C(_136_), .Y(_137_) );
NOR2X1 NOR2X1_19 ( .A(_134_), .B(_137_), .Y(_138_) );
NAND2X1 NAND2X1_20 ( .A(asr1_rom_3__4_), .B(_34_), .Y(_139_) );
NAND3X1 NAND3X1_33 ( .A(asr1_rom_4__4_), .B(_36__bF_buf3), .C(_4__bF_buf1), .Y(_140_) );
NAND3X1 NAND3X1_34 ( .A(asr1_rom_0__4_), .B(_20_), .C(_36__bF_buf2), .Y(_141_) );
NAND3X1 NAND3X1_35 ( .A(asr1_en_4_), .B(_29_), .C(_33__bF_buf2), .Y(_142_) );
AND2X2 AND2X2_10 ( .A(_142_), .B(_141_), .Y(_143_) );
NAND3X1 NAND3X1_36 ( .A(_139_), .B(_140_), .C(_143_), .Y(_144_) );
NAND3X1 NAND3X1_37 ( .A(asr1_rom_7__4_), .B(_33__bF_buf1), .C(_4__bF_buf0), .Y(_145_) );
NAND3X1 NAND3X1_38 ( .A(asr1_rom_8__4_), .B(_36__bF_buf1), .C(_13_), .Y(_146_) );
AOI22X1 AOI22X1_5 ( .A(_46_), .B(asr1_rom_12__4_), .C(asr1_rom_11__4_), .D(_45_), .Y(_147_) );
NAND3X1 NAND3X1_39 ( .A(_145_), .B(_146_), .C(_147_), .Y(_148_) );
NOR2X1 NOR2X1_20 ( .A(_144_), .B(_148_), .Y(_149_) );
NAND3X1 NAND3X1_40 ( .A(_131_), .B(_138_), .C(_149_), .Y(asr1_dataout_4_) );
INVX1 INVX1_38 ( .A(asr1_rom_6__5_), .Y(_150_) );
INVX1 INVX1_39 ( .A(asr1_rom_5__5_), .Y(_151_) );
OAI22X1 OAI22X1_16 ( .A(_150_), .B(_9_), .C(_151_), .D(_7_), .Y(_152_) );
INVX1 INVX1_40 ( .A(asr1_rom_10__5_), .Y(_153_) );
INVX1 INVX1_41 ( .A(asr1_rom_9__5_), .Y(_154_) );
OAI22X1 OAI22X1_17 ( .A(_153_), .B(_15_), .C(_154_), .D(_14_), .Y(_155_) );
NOR2X1 NOR2X1_21 ( .A(_155_), .B(_152_), .Y(_156_) );
INVX1 INVX1_42 ( .A(asr1_rom_2__5_), .Y(_157_) );
INVX1 INVX1_43 ( .A(asr1_rom_1__5_), .Y(_158_) );
OAI22X1 OAI22X1_18 ( .A(_157_), .B(_22_), .C(_158_), .D(_21_), .Y(_159_) );
INVX1 INVX1_44 ( .A(asr1_rom_14__5_), .Y(_160_) );
NAND2X1 NAND2X1_21 ( .A(asr1_rom_13__5_), .B(_27_), .Y(_161_) );
OAI21X1 OAI21X1_6 ( .A(_160_), .B(_30_), .C(_161_), .Y(_162_) );
NOR2X1 NOR2X1_22 ( .A(_159_), .B(_162_), .Y(_163_) );
NAND2X1 NAND2X1_22 ( .A(asr1_rom_3__5_), .B(_34_), .Y(_164_) );
NAND3X1 NAND3X1_41 ( .A(asr1_rom_4__5_), .B(_36__bF_buf0), .C(_4__bF_buf3), .Y(_165_) );
NAND3X1 NAND3X1_42 ( .A(asr1_rom_0__5_), .B(_20_), .C(_36__bF_buf3), .Y(_166_) );
NAND3X1 NAND3X1_43 ( .A(asr1_en_5_), .B(_29_), .C(_33__bF_buf0), .Y(_167_) );
AND2X2 AND2X2_11 ( .A(_167_), .B(_166_), .Y(_168_) );
NAND3X1 NAND3X1_44 ( .A(_164_), .B(_165_), .C(_168_), .Y(_169_) );
NAND3X1 NAND3X1_45 ( .A(asr1_rom_7__5_), .B(_33__bF_buf3), .C(_4__bF_buf2), .Y(_170_) );
NAND3X1 NAND3X1_46 ( .A(asr1_rom_8__5_), .B(_36__bF_buf2), .C(_13_), .Y(_171_) );
AOI22X1 AOI22X1_6 ( .A(_46_), .B(asr1_rom_12__5_), .C(asr1_rom_11__5_), .D(_45_), .Y(_172_) );
NAND3X1 NAND3X1_47 ( .A(_170_), .B(_171_), .C(_172_), .Y(_173_) );
NOR2X1 NOR2X1_23 ( .A(_169_), .B(_173_), .Y(_174_) );
NAND3X1 NAND3X1_48 ( .A(_156_), .B(_163_), .C(_174_), .Y(asr1_dataout_5_) );
INVX1 INVX1_45 ( .A(asr1_rom_6__6_), .Y(_175_) );
INVX1 INVX1_46 ( .A(asr1_rom_5__6_), .Y(_176_) );
OAI22X1 OAI22X1_19 ( .A(_175_), .B(_9_), .C(_176_), .D(_7_), .Y(_177_) );
INVX1 INVX1_47 ( .A(asr1_rom_10__6_), .Y(_178_) );
INVX1 INVX1_48 ( .A(asr1_rom_9__6_), .Y(_179_) );
OAI22X1 OAI22X1_20 ( .A(_178_), .B(_15_), .C(_179_), .D(_14_), .Y(_180_) );
NOR2X1 NOR2X1_24 ( .A(_180_), .B(_177_), .Y(_181_) );
INVX1 INVX1_49 ( .A(asr1_rom_2__6_), .Y(_182_) );
INVX1 INVX1_50 ( .A(asr1_rom_1__6_), .Y(_183_) );
OAI22X1 OAI22X1_21 ( .A(_182_), .B(_22_), .C(_183_), .D(_21_), .Y(_184_) );
INVX1 INVX1_51 ( .A(asr1_rom_14__6_), .Y(_185_) );
NAND2X1 NAND2X1_23 ( .A(asr1_rom_13__6_), .B(_27_), .Y(_186_) );
OAI21X1 OAI21X1_7 ( .A(_185_), .B(_30_), .C(_186_), .Y(_187_) );
NOR2X1 NOR2X1_25 ( .A(_184_), .B(_187_), .Y(_188_) );
NAND2X1 NAND2X1_24 ( .A(asr1_rom_3__6_), .B(_34_), .Y(_189_) );
NAND3X1 NAND3X1_49 ( .A(asr1_rom_4__6_), .B(_36__bF_buf1), .C(_4__bF_buf1), .Y(_190_) );
NAND3X1 NAND3X1_50 ( .A(asr1_rom_0__6_), .B(_20_), .C(_36__bF_buf0), .Y(_191_) );
NAND3X1 NAND3X1_51 ( .A(asr1_en_6_), .B(_29_), .C(_33__bF_buf2), .Y(_192_) );
AND2X2 AND2X2_12 ( .A(_192_), .B(_191_), .Y(_193_) );
NAND3X1 NAND3X1_52 ( .A(_189_), .B(_190_), .C(_193_), .Y(_194_) );
NAND3X1 NAND3X1_53 ( .A(asr1_rom_7__6_), .B(_33__bF_buf1), .C(_4__bF_buf0), .Y(_195_) );
NAND3X1 NAND3X1_54 ( .A(asr1_rom_8__6_), .B(_36__bF_buf3), .C(_13_), .Y(_196_) );
AOI22X1 AOI22X1_7 ( .A(_46_), .B(asr1_rom_12__6_), .C(asr1_rom_11__6_), .D(_45_), .Y(_197_) );
NAND3X1 NAND3X1_55 ( .A(_195_), .B(_196_), .C(_197_), .Y(_198_) );
NOR2X1 NOR2X1_26 ( .A(_194_), .B(_198_), .Y(_199_) );
NAND3X1 NAND3X1_56 ( .A(_181_), .B(_188_), .C(_199_), .Y(asr1_dataout_6_) );
INVX1 INVX1_52 ( .A(asr1_rom_6__7_), .Y(_200_) );
INVX1 INVX1_53 ( .A(asr1_rom_5__7_), .Y(_201_) );
OAI22X1 OAI22X1_22 ( .A(_200_), .B(_9_), .C(_201_), .D(_7_), .Y(_202_) );
INVX1 INVX1_54 ( .A(asr1_rom_10__7_), .Y(_203_) );
INVX1 INVX1_55 ( .A(asr1_rom_9__7_), .Y(_204_) );
OAI22X1 OAI22X1_23 ( .A(_203_), .B(_15_), .C(_204_), .D(_14_), .Y(_205_) );
NOR2X1 NOR2X1_27 ( .A(_205_), .B(_202_), .Y(_206_) );
INVX1 INVX1_56 ( .A(asr1_rom_2__7_), .Y(_207_) );
INVX1 INVX1_57 ( .A(asr1_rom_1__7_), .Y(_208_) );
OAI22X1 OAI22X1_24 ( .A(_207_), .B(_22_), .C(_208_), .D(_21_), .Y(_209_) );
INVX1 INVX1_58 ( .A(asr1_rom_14__7_), .Y(_210_) );
NAND2X1 NAND2X1_25 ( .A(asr1_rom_13__7_), .B(_27_), .Y(_211_) );
OAI21X1 OAI21X1_8 ( .A(_210_), .B(_30_), .C(_211_), .Y(_212_) );
NOR2X1 NOR2X1_28 ( .A(_209_), .B(_212_), .Y(_213_) );
NAND2X1 NAND2X1_26 ( .A(asr1_rom_3__7_), .B(_34_), .Y(_214_) );
NAND3X1 NAND3X1_57 ( .A(asr1_rom_4__7_), .B(_36__bF_buf2), .C(_4__bF_buf3), .Y(_215_) );
NAND3X1 NAND3X1_58 ( .A(asr1_rom_0__7_), .B(_20_), .C(_36__bF_buf1), .Y(_216_) );
NAND3X1 NAND3X1_59 ( .A(asr1_en_7_), .B(_29_), .C(_33__bF_buf0), .Y(_217_) );
AND2X2 AND2X2_13 ( .A(_217_), .B(_216_), .Y(_218_) );
NAND3X1 NAND3X1_60 ( .A(_214_), .B(_215_), .C(_218_), .Y(_219_) );
NAND3X1 NAND3X1_61 ( .A(asr1_rom_7__7_), .B(_33__bF_buf3), .C(_4__bF_buf2), .Y(_220_) );
NAND3X1 NAND3X1_62 ( .A(asr1_rom_8__7_), .B(_36__bF_buf0), .C(_13_), .Y(_221_) );
AOI22X1 AOI22X1_8 ( .A(_46_), .B(asr1_rom_12__7_), .C(asr1_rom_11__7_), .D(_45_), .Y(_222_) );
NAND3X1 NAND3X1_63 ( .A(_220_), .B(_221_), .C(_222_), .Y(_223_) );
NOR2X1 NOR2X1_29 ( .A(_219_), .B(_223_), .Y(_224_) );
NAND3X1 NAND3X1_64 ( .A(_206_), .B(_213_), .C(_224_), .Y(asr1_dataout_7_) );
INVX1 INVX1_59 ( .A(rst_bF_buf5), .Y(_0_) );
DFFSR DFFSR_1 ( .CLK(clk2_clkout_bF_buf41), .D(reg1_dataout_0_), .Q(asr1_rom_0__0_), .R(_0__bF_buf10), .S(vdd) );
DFFSR DFFSR_2 ( .CLK(clk2_clkout_bF_buf40), .D(reg1_dataout_1_), .Q(asr1_rom_0__1_), .R(_0__bF_buf9), .S(vdd) );
DFFSR DFFSR_3 ( .CLK(clk2_clkout_bF_buf39), .D(reg1_dataout_2_), .Q(asr1_rom_0__2_), .R(_0__bF_buf8), .S(vdd) );
DFFSR DFFSR_4 ( .CLK(clk2_clkout_bF_buf38), .D(reg1_dataout_3_), .Q(asr1_rom_0__3_), .R(_0__bF_buf7), .S(vdd) );
DFFSR DFFSR_5 ( .CLK(clk2_clkout_bF_buf37), .D(reg1_dataout_4_), .Q(asr1_rom_0__4_), .R(_0__bF_buf6), .S(vdd) );
DFFSR DFFSR_6 ( .CLK(clk2_clkout_bF_buf36), .D(reg1_dataout_5_), .Q(asr1_rom_0__5_), .R(_0__bF_buf5), .S(vdd) );
DFFSR DFFSR_7 ( .CLK(clk2_clkout_bF_buf35), .D(reg1_dataout_6_), .Q(asr1_rom_0__6_), .R(_0__bF_buf4), .S(vdd) );
DFFSR DFFSR_8 ( .CLK(clk2_clkout_bF_buf34), .D(reg1_dataout_7_), .Q(asr1_rom_0__7_), .R(_0__bF_buf3), .S(vdd) );
DFFSR DFFSR_9 ( .CLK(clk2_clkout_bF_buf33), .D(asr1_rom_6__0_), .Q(asr1_rom_7__0_), .R(_0__bF_buf2), .S(vdd) );
DFFSR DFFSR_10 ( .CLK(clk2_clkout_bF_buf32), .D(asr1_rom_6__1_), .Q(asr1_rom_7__1_), .R(_0__bF_buf1), .S(vdd) );
DFFSR DFFSR_11 ( .CLK(clk2_clkout_bF_buf31), .D(asr1_rom_6__2_), .Q(asr1_rom_7__2_), .R(_0__bF_buf0), .S(vdd) );
DFFSR DFFSR_12 ( .CLK(clk2_clkout_bF_buf30), .D(asr1_rom_6__3_), .Q(asr1_rom_7__3_), .R(_0__bF_buf10), .S(vdd) );
DFFSR DFFSR_13 ( .CLK(clk2_clkout_bF_buf29), .D(asr1_rom_6__4_), .Q(asr1_rom_7__4_), .R(_0__bF_buf9), .S(vdd) );
DFFSR DFFSR_14 ( .CLK(clk2_clkout_bF_buf28), .D(asr1_rom_6__5_), .Q(asr1_rom_7__5_), .R(_0__bF_buf8), .S(vdd) );
DFFSR DFFSR_15 ( .CLK(clk2_clkout_bF_buf27), .D(asr1_rom_6__6_), .Q(asr1_rom_7__6_), .R(_0__bF_buf7), .S(vdd) );
DFFSR DFFSR_16 ( .CLK(clk2_clkout_bF_buf26), .D(asr1_rom_6__7_), .Q(asr1_rom_7__7_), .R(_0__bF_buf6), .S(vdd) );
DFFSR DFFSR_17 ( .CLK(clk2_clkout_bF_buf25), .D(asr1_rom_1__0_), .Q(asr1_rom_2__0_), .R(_0__bF_buf5), .S(vdd) );
DFFSR DFFSR_18 ( .CLK(clk2_clkout_bF_buf24), .D(asr1_rom_1__1_), .Q(asr1_rom_2__1_), .R(_0__bF_buf4), .S(vdd) );
DFFSR DFFSR_19 ( .CLK(clk2_clkout_bF_buf23), .D(asr1_rom_1__2_), .Q(asr1_rom_2__2_), .R(_0__bF_buf3), .S(vdd) );
DFFSR DFFSR_20 ( .CLK(clk2_clkout_bF_buf22), .D(asr1_rom_1__3_), .Q(asr1_rom_2__3_), .R(_0__bF_buf2), .S(vdd) );
DFFSR DFFSR_21 ( .CLK(clk2_clkout_bF_buf21), .D(asr1_rom_1__4_), .Q(asr1_rom_2__4_), .R(_0__bF_buf1), .S(vdd) );
DFFSR DFFSR_22 ( .CLK(clk2_clkout_bF_buf20), .D(asr1_rom_1__5_), .Q(asr1_rom_2__5_), .R(_0__bF_buf0), .S(vdd) );
DFFSR DFFSR_23 ( .CLK(clk2_clkout_bF_buf19), .D(asr1_rom_1__6_), .Q(asr1_rom_2__6_), .R(_0__bF_buf10), .S(vdd) );
DFFSR DFFSR_24 ( .CLK(clk2_clkout_bF_buf18), .D(asr1_rom_1__7_), .Q(asr1_rom_2__7_), .R(_0__bF_buf9), .S(vdd) );
DFFSR DFFSR_25 ( .CLK(clk2_clkout_bF_buf17), .D(asr1_rom_0__0_), .Q(asr1_rom_1__0_), .R(_0__bF_buf8), .S(vdd) );
DFFSR DFFSR_26 ( .CLK(clk2_clkout_bF_buf16), .D(asr1_rom_0__1_), .Q(asr1_rom_1__1_), .R(_0__bF_buf7), .S(vdd) );
DFFSR DFFSR_27 ( .CLK(clk2_clkout_bF_buf15), .D(asr1_rom_0__2_), .Q(asr1_rom_1__2_), .R(_0__bF_buf6), .S(vdd) );
DFFSR DFFSR_28 ( .CLK(clk2_clkout_bF_buf14), .D(asr1_rom_0__3_), .Q(asr1_rom_1__3_), .R(_0__bF_buf5), .S(vdd) );
DFFSR DFFSR_29 ( .CLK(clk2_clkout_bF_buf13), .D(asr1_rom_0__4_), .Q(asr1_rom_1__4_), .R(_0__bF_buf4), .S(vdd) );
DFFSR DFFSR_30 ( .CLK(clk2_clkout_bF_buf12), .D(asr1_rom_0__5_), .Q(asr1_rom_1__5_), .R(_0__bF_buf3), .S(vdd) );
DFFSR DFFSR_31 ( .CLK(clk2_clkout_bF_buf11), .D(asr1_rom_0__6_), .Q(asr1_rom_1__6_), .R(_0__bF_buf2), .S(vdd) );
DFFSR DFFSR_32 ( .CLK(clk2_clkout_bF_buf10), .D(asr1_rom_0__7_), .Q(asr1_rom_1__7_), .R(_0__bF_buf1), .S(vdd) );
DFFSR DFFSR_33 ( .CLK(clk2_clkout_bF_buf9), .D(asr1_rom_2__0_), .Q(asr1_rom_3__0_), .R(_0__bF_buf0), .S(vdd) );
DFFSR DFFSR_34 ( .CLK(clk2_clkout_bF_buf8), .D(asr1_rom_2__1_), .Q(asr1_rom_3__1_), .R(_0__bF_buf10), .S(vdd) );
DFFSR DFFSR_35 ( .CLK(clk2_clkout_bF_buf7), .D(asr1_rom_2__2_), .Q(asr1_rom_3__2_), .R(_0__bF_buf9), .S(vdd) );
DFFSR DFFSR_36 ( .CLK(clk2_clkout_bF_buf6), .D(asr1_rom_2__3_), .Q(asr1_rom_3__3_), .R(_0__bF_buf8), .S(vdd) );
DFFSR DFFSR_37 ( .CLK(clk2_clkout_bF_buf5), .D(asr1_rom_2__4_), .Q(asr1_rom_3__4_), .R(_0__bF_buf7), .S(vdd) );
DFFSR DFFSR_38 ( .CLK(clk2_clkout_bF_buf4), .D(asr1_rom_2__5_), .Q(asr1_rom_3__5_), .R(_0__bF_buf6), .S(vdd) );
DFFSR DFFSR_39 ( .CLK(clk2_clkout_bF_buf3), .D(asr1_rom_2__6_), .Q(asr1_rom_3__6_), .R(_0__bF_buf5), .S(vdd) );
DFFSR DFFSR_40 ( .CLK(clk2_clkout_bF_buf2), .D(asr1_rom_2__7_), .Q(asr1_rom_3__7_), .R(_0__bF_buf4), .S(vdd) );
DFFSR DFFSR_41 ( .CLK(clk2_clkout_bF_buf1), .D(asr1_rom_3__0_), .Q(asr1_rom_4__0_), .R(_0__bF_buf3), .S(vdd) );
DFFSR DFFSR_42 ( .CLK(clk2_clkout_bF_buf0), .D(asr1_rom_3__1_), .Q(asr1_rom_4__1_), .R(_0__bF_buf2), .S(vdd) );
DFFSR DFFSR_43 ( .CLK(clk2_clkout_bF_buf41), .D(asr1_rom_3__2_), .Q(asr1_rom_4__2_), .R(_0__bF_buf1), .S(vdd) );
DFFSR DFFSR_44 ( .CLK(clk2_clkout_bF_buf40), .D(asr1_rom_3__3_), .Q(asr1_rom_4__3_), .R(_0__bF_buf0), .S(vdd) );
DFFSR DFFSR_45 ( .CLK(clk2_clkout_bF_buf39), .D(asr1_rom_3__4_), .Q(asr1_rom_4__4_), .R(_0__bF_buf10), .S(vdd) );
DFFSR DFFSR_46 ( .CLK(clk2_clkout_bF_buf38), .D(asr1_rom_3__5_), .Q(asr1_rom_4__5_), .R(_0__bF_buf9), .S(vdd) );
DFFSR DFFSR_47 ( .CLK(clk2_clkout_bF_buf37), .D(asr1_rom_3__6_), .Q(asr1_rom_4__6_), .R(_0__bF_buf8), .S(vdd) );
DFFSR DFFSR_48 ( .CLK(clk2_clkout_bF_buf36), .D(asr1_rom_3__7_), .Q(asr1_rom_4__7_), .R(_0__bF_buf7), .S(vdd) );
DFFSR DFFSR_49 ( .CLK(clk2_clkout_bF_buf35), .D(asr1_rom_5__0_), .Q(asr1_rom_6__0_), .R(_0__bF_buf6), .S(vdd) );
DFFSR DFFSR_50 ( .CLK(clk2_clkout_bF_buf34), .D(asr1_rom_5__1_), .Q(asr1_rom_6__1_), .R(_0__bF_buf5), .S(vdd) );
DFFSR DFFSR_51 ( .CLK(clk2_clkout_bF_buf33), .D(asr1_rom_5__2_), .Q(asr1_rom_6__2_), .R(_0__bF_buf4), .S(vdd) );
DFFSR DFFSR_52 ( .CLK(clk2_clkout_bF_buf32), .D(asr1_rom_5__3_), .Q(asr1_rom_6__3_), .R(_0__bF_buf3), .S(vdd) );
DFFSR DFFSR_53 ( .CLK(clk2_clkout_bF_buf31), .D(asr1_rom_5__4_), .Q(asr1_rom_6__4_), .R(_0__bF_buf2), .S(vdd) );
DFFSR DFFSR_54 ( .CLK(clk2_clkout_bF_buf30), .D(asr1_rom_5__5_), .Q(asr1_rom_6__5_), .R(_0__bF_buf1), .S(vdd) );
DFFSR DFFSR_55 ( .CLK(clk2_clkout_bF_buf29), .D(asr1_rom_5__6_), .Q(asr1_rom_6__6_), .R(_0__bF_buf0), .S(vdd) );
DFFSR DFFSR_56 ( .CLK(clk2_clkout_bF_buf28), .D(asr1_rom_5__7_), .Q(asr1_rom_6__7_), .R(_0__bF_buf10), .S(vdd) );
DFFSR DFFSR_57 ( .CLK(clk2_clkout_bF_buf27), .D(asr1_rom_4__0_), .Q(asr1_rom_5__0_), .R(_0__bF_buf9), .S(vdd) );
DFFSR DFFSR_58 ( .CLK(clk2_clkout_bF_buf26), .D(asr1_rom_4__1_), .Q(asr1_rom_5__1_), .R(_0__bF_buf8), .S(vdd) );
DFFSR DFFSR_59 ( .CLK(clk2_clkout_bF_buf25), .D(asr1_rom_4__2_), .Q(asr1_rom_5__2_), .R(_0__bF_buf7), .S(vdd) );
DFFSR DFFSR_60 ( .CLK(clk2_clkout_bF_buf24), .D(asr1_rom_4__3_), .Q(asr1_rom_5__3_), .R(_0__bF_buf6), .S(vdd) );
DFFSR DFFSR_61 ( .CLK(clk2_clkout_bF_buf23), .D(asr1_rom_4__4_), .Q(asr1_rom_5__4_), .R(_0__bF_buf5), .S(vdd) );
DFFSR DFFSR_62 ( .CLK(clk2_clkout_bF_buf22), .D(asr1_rom_4__5_), .Q(asr1_rom_5__5_), .R(_0__bF_buf4), .S(vdd) );
DFFSR DFFSR_63 ( .CLK(clk2_clkout_bF_buf21), .D(asr1_rom_4__6_), .Q(asr1_rom_5__6_), .R(_0__bF_buf3), .S(vdd) );
DFFSR DFFSR_64 ( .CLK(clk2_clkout_bF_buf20), .D(asr1_rom_4__7_), .Q(asr1_rom_5__7_), .R(_0__bF_buf2), .S(vdd) );
DFFSR DFFSR_65 ( .CLK(clk2_clkout_bF_buf19), .D(asr1_rom_7__0_), .Q(asr1_rom_8__0_), .R(_0__bF_buf1), .S(vdd) );
DFFSR DFFSR_66 ( .CLK(clk2_clkout_bF_buf18), .D(asr1_rom_7__1_), .Q(asr1_rom_8__1_), .R(_0__bF_buf0), .S(vdd) );
DFFSR DFFSR_67 ( .CLK(clk2_clkout_bF_buf17), .D(asr1_rom_7__2_), .Q(asr1_rom_8__2_), .R(_0__bF_buf10), .S(vdd) );
DFFSR DFFSR_68 ( .CLK(clk2_clkout_bF_buf16), .D(asr1_rom_7__3_), .Q(asr1_rom_8__3_), .R(_0__bF_buf9), .S(vdd) );
DFFSR DFFSR_69 ( .CLK(clk2_clkout_bF_buf15), .D(asr1_rom_7__4_), .Q(asr1_rom_8__4_), .R(_0__bF_buf8), .S(vdd) );
DFFSR DFFSR_70 ( .CLK(clk2_clkout_bF_buf14), .D(asr1_rom_7__5_), .Q(asr1_rom_8__5_), .R(_0__bF_buf7), .S(vdd) );
DFFSR DFFSR_71 ( .CLK(clk2_clkout_bF_buf13), .D(asr1_rom_7__6_), .Q(asr1_rom_8__6_), .R(_0__bF_buf6), .S(vdd) );
DFFSR DFFSR_72 ( .CLK(clk2_clkout_bF_buf12), .D(asr1_rom_7__7_), .Q(asr1_rom_8__7_), .R(_0__bF_buf5), .S(vdd) );
DFFSR DFFSR_73 ( .CLK(clk2_clkout_bF_buf11), .D(asr1_rom_8__0_), .Q(asr1_rom_9__0_), .R(_0__bF_buf4), .S(vdd) );
DFFSR DFFSR_74 ( .CLK(clk2_clkout_bF_buf10), .D(asr1_rom_8__1_), .Q(asr1_rom_9__1_), .R(_0__bF_buf3), .S(vdd) );
DFFSR DFFSR_75 ( .CLK(clk2_clkout_bF_buf9), .D(asr1_rom_8__2_), .Q(asr1_rom_9__2_), .R(_0__bF_buf2), .S(vdd) );
DFFSR DFFSR_76 ( .CLK(clk2_clkout_bF_buf8), .D(asr1_rom_8__3_), .Q(asr1_rom_9__3_), .R(_0__bF_buf1), .S(vdd) );
DFFSR DFFSR_77 ( .CLK(clk2_clkout_bF_buf7), .D(asr1_rom_8__4_), .Q(asr1_rom_9__4_), .R(_0__bF_buf0), .S(vdd) );
DFFSR DFFSR_78 ( .CLK(clk2_clkout_bF_buf6), .D(asr1_rom_8__5_), .Q(asr1_rom_9__5_), .R(_0__bF_buf10), .S(vdd) );
DFFSR DFFSR_79 ( .CLK(clk2_clkout_bF_buf5), .D(asr1_rom_8__6_), .Q(asr1_rom_9__6_), .R(_0__bF_buf9), .S(vdd) );
DFFSR DFFSR_80 ( .CLK(clk2_clkout_bF_buf4), .D(asr1_rom_8__7_), .Q(asr1_rom_9__7_), .R(_0__bF_buf8), .S(vdd) );
DFFSR DFFSR_81 ( .CLK(clk2_clkout_bF_buf3), .D(asr1_rom_9__0_), .Q(asr1_rom_10__0_), .R(_0__bF_buf7), .S(vdd) );
DFFSR DFFSR_82 ( .CLK(clk2_clkout_bF_buf2), .D(asr1_rom_9__1_), .Q(asr1_rom_10__1_), .R(_0__bF_buf6), .S(vdd) );
DFFSR DFFSR_83 ( .CLK(clk2_clkout_bF_buf1), .D(asr1_rom_9__2_), .Q(asr1_rom_10__2_), .R(_0__bF_buf5), .S(vdd) );
DFFSR DFFSR_84 ( .CLK(clk2_clkout_bF_buf0), .D(asr1_rom_9__3_), .Q(asr1_rom_10__3_), .R(_0__bF_buf4), .S(vdd) );
DFFSR DFFSR_85 ( .CLK(clk2_clkout_bF_buf41), .D(asr1_rom_9__4_), .Q(asr1_rom_10__4_), .R(_0__bF_buf3), .S(vdd) );
DFFSR DFFSR_86 ( .CLK(clk2_clkout_bF_buf40), .D(asr1_rom_9__5_), .Q(asr1_rom_10__5_), .R(_0__bF_buf2), .S(vdd) );
DFFSR DFFSR_87 ( .CLK(clk2_clkout_bF_buf39), .D(asr1_rom_9__6_), .Q(asr1_rom_10__6_), .R(_0__bF_buf1), .S(vdd) );
DFFSR DFFSR_88 ( .CLK(clk2_clkout_bF_buf38), .D(asr1_rom_9__7_), .Q(asr1_rom_10__7_), .R(_0__bF_buf0), .S(vdd) );
DFFSR DFFSR_89 ( .CLK(clk2_clkout_bF_buf37), .D(asr1_rom_10__0_), .Q(asr1_rom_11__0_), .R(_0__bF_buf10), .S(vdd) );
DFFSR DFFSR_90 ( .CLK(clk2_clkout_bF_buf36), .D(asr1_rom_10__1_), .Q(asr1_rom_11__1_), .R(_0__bF_buf9), .S(vdd) );
DFFSR DFFSR_91 ( .CLK(clk2_clkout_bF_buf35), .D(asr1_rom_10__2_), .Q(asr1_rom_11__2_), .R(_0__bF_buf8), .S(vdd) );
DFFSR DFFSR_92 ( .CLK(clk2_clkout_bF_buf34), .D(asr1_rom_10__3_), .Q(asr1_rom_11__3_), .R(_0__bF_buf7), .S(vdd) );
DFFSR DFFSR_93 ( .CLK(clk2_clkout_bF_buf33), .D(asr1_rom_10__4_), .Q(asr1_rom_11__4_), .R(_0__bF_buf6), .S(vdd) );
DFFSR DFFSR_94 ( .CLK(clk2_clkout_bF_buf32), .D(asr1_rom_10__5_), .Q(asr1_rom_11__5_), .R(_0__bF_buf5), .S(vdd) );
DFFSR DFFSR_95 ( .CLK(clk2_clkout_bF_buf31), .D(asr1_rom_10__6_), .Q(asr1_rom_11__6_), .R(_0__bF_buf4), .S(vdd) );
DFFSR DFFSR_96 ( .CLK(clk2_clkout_bF_buf30), .D(asr1_rom_10__7_), .Q(asr1_rom_11__7_), .R(_0__bF_buf3), .S(vdd) );
DFFSR DFFSR_97 ( .CLK(clk2_clkout_bF_buf29), .D(asr1_rom_11__0_), .Q(asr1_rom_12__0_), .R(_0__bF_buf2), .S(vdd) );
DFFSR DFFSR_98 ( .CLK(clk2_clkout_bF_buf28), .D(asr1_rom_11__1_), .Q(asr1_rom_12__1_), .R(_0__bF_buf1), .S(vdd) );
DFFSR DFFSR_99 ( .CLK(clk2_clkout_bF_buf27), .D(asr1_rom_11__2_), .Q(asr1_rom_12__2_), .R(_0__bF_buf0), .S(vdd) );
DFFSR DFFSR_100 ( .CLK(clk2_clkout_bF_buf26), .D(asr1_rom_11__3_), .Q(asr1_rom_12__3_), .R(_0__bF_buf10), .S(vdd) );
DFFSR DFFSR_101 ( .CLK(clk2_clkout_bF_buf25), .D(asr1_rom_11__4_), .Q(asr1_rom_12__4_), .R(_0__bF_buf9), .S(vdd) );
DFFSR DFFSR_102 ( .CLK(clk2_clkout_bF_buf24), .D(asr1_rom_11__5_), .Q(asr1_rom_12__5_), .R(_0__bF_buf8), .S(vdd) );
DFFSR DFFSR_103 ( .CLK(clk2_clkout_bF_buf23), .D(asr1_rom_11__6_), .Q(asr1_rom_12__6_), .R(_0__bF_buf7), .S(vdd) );
DFFSR DFFSR_104 ( .CLK(clk2_clkout_bF_buf22), .D(asr1_rom_11__7_), .Q(asr1_rom_12__7_), .R(_0__bF_buf6), .S(vdd) );
DFFSR DFFSR_105 ( .CLK(clk2_clkout_bF_buf21), .D(asr1_rom_12__0_), .Q(asr1_rom_13__0_), .R(_0__bF_buf5), .S(vdd) );
DFFSR DFFSR_106 ( .CLK(clk2_clkout_bF_buf20), .D(asr1_rom_12__1_), .Q(asr1_rom_13__1_), .R(_0__bF_buf4), .S(vdd) );
DFFSR DFFSR_107 ( .CLK(clk2_clkout_bF_buf19), .D(asr1_rom_12__2_), .Q(asr1_rom_13__2_), .R(_0__bF_buf3), .S(vdd) );
DFFSR DFFSR_108 ( .CLK(clk2_clkout_bF_buf18), .D(asr1_rom_12__3_), .Q(asr1_rom_13__3_), .R(_0__bF_buf2), .S(vdd) );
DFFSR DFFSR_109 ( .CLK(clk2_clkout_bF_buf17), .D(asr1_rom_12__4_), .Q(asr1_rom_13__4_), .R(_0__bF_buf1), .S(vdd) );
DFFSR DFFSR_110 ( .CLK(clk2_clkout_bF_buf16), .D(asr1_rom_12__5_), .Q(asr1_rom_13__5_), .R(_0__bF_buf0), .S(vdd) );
DFFSR DFFSR_111 ( .CLK(clk2_clkout_bF_buf15), .D(asr1_rom_12__6_), .Q(asr1_rom_13__6_), .R(_0__bF_buf10), .S(vdd) );
DFFSR DFFSR_112 ( .CLK(clk2_clkout_bF_buf14), .D(asr1_rom_12__7_), .Q(asr1_rom_13__7_), .R(_0__bF_buf9), .S(vdd) );
DFFSR DFFSR_113 ( .CLK(clk2_clkout_bF_buf13), .D(asr1_rom_13__0_), .Q(asr1_rom_14__0_), .R(_0__bF_buf8), .S(vdd) );
DFFSR DFFSR_114 ( .CLK(clk2_clkout_bF_buf12), .D(asr1_rom_13__1_), .Q(asr1_rom_14__1_), .R(_0__bF_buf7), .S(vdd) );
DFFSR DFFSR_115 ( .CLK(clk2_clkout_bF_buf11), .D(asr1_rom_13__2_), .Q(asr1_rom_14__2_), .R(_0__bF_buf6), .S(vdd) );
DFFSR DFFSR_116 ( .CLK(clk2_clkout_bF_buf10), .D(asr1_rom_13__3_), .Q(asr1_rom_14__3_), .R(_0__bF_buf5), .S(vdd) );
DFFSR DFFSR_117 ( .CLK(clk2_clkout_bF_buf9), .D(asr1_rom_13__4_), .Q(asr1_rom_14__4_), .R(_0__bF_buf4), .S(vdd) );
DFFSR DFFSR_118 ( .CLK(clk2_clkout_bF_buf8), .D(asr1_rom_13__5_), .Q(asr1_rom_14__5_), .R(_0__bF_buf3), .S(vdd) );
DFFSR DFFSR_119 ( .CLK(clk2_clkout_bF_buf7), .D(asr1_rom_13__6_), .Q(asr1_rom_14__6_), .R(_0__bF_buf2), .S(vdd) );
DFFSR DFFSR_120 ( .CLK(clk2_clkout_bF_buf6), .D(asr1_rom_13__7_), .Q(asr1_rom_14__7_), .R(_0__bF_buf1), .S(vdd) );
DFFSR DFFSR_121 ( .CLK(clk2_clkout_bF_buf5), .D(asr1_rom_14__0_), .Q(asr1_en_0_), .R(_0__bF_buf0), .S(vdd) );
DFFSR DFFSR_122 ( .CLK(clk2_clkout_bF_buf4), .D(asr1_rom_14__1_), .Q(asr1_en_1_), .R(_0__bF_buf10), .S(vdd) );
DFFSR DFFSR_123 ( .CLK(clk2_clkout_bF_buf3), .D(asr1_rom_14__2_), .Q(asr1_en_2_), .R(_0__bF_buf9), .S(vdd) );
DFFSR DFFSR_124 ( .CLK(clk2_clkout_bF_buf2), .D(asr1_rom_14__3_), .Q(asr1_en_3_), .R(_0__bF_buf8), .S(vdd) );
DFFSR DFFSR_125 ( .CLK(clk2_clkout_bF_buf1), .D(asr1_rom_14__4_), .Q(asr1_en_4_), .R(_0__bF_buf7), .S(vdd) );
DFFSR DFFSR_126 ( .CLK(clk2_clkout_bF_buf0), .D(asr1_rom_14__5_), .Q(asr1_en_5_), .R(_0__bF_buf6), .S(vdd) );
DFFSR DFFSR_127 ( .CLK(clk2_clkout_bF_buf41), .D(asr1_rom_14__6_), .Q(asr1_en_6_), .R(_0__bF_buf5), .S(vdd) );
DFFSR DFFSR_128 ( .CLK(clk2_clkout_bF_buf40), .D(asr1_rom_14__7_), .Q(asr1_en_7_), .R(_0__bF_buf4), .S(vdd) );
INVX1 INVX1_60 ( .A(asr2_rom_6__0_), .Y(_226_) );
INVX1 INVX1_61 ( .A(asr2_rom_5__0_), .Y(_227_) );
INVX1 INVX1_62 ( .A(counterdown_counter_3_), .Y(_228_) );
AND2X2 AND2X2_14 ( .A(_228_), .B(counterdown_counter_2_), .Y(_229_) );
INVX1 INVX1_63 ( .A(counterdown_counter_1_), .Y(_230_) );
AND2X2 AND2X2_15 ( .A(_230_), .B(counterdown_counter_0_), .Y(_231_) );
NAND2X1 NAND2X1_27 ( .A(_229__bF_buf3), .B(_231_), .Y(_232_) );
NOR2X1 NOR2X1_30 ( .A(counterdown_counter_0_), .B(_230_), .Y(_233_) );
NAND2X1 NAND2X1_28 ( .A(_233_), .B(_229__bF_buf2), .Y(_234_) );
OAI22X1 OAI22X1_25 ( .A(_226_), .B(_234_), .C(_227_), .D(_232_), .Y(_235_) );
INVX1 INVX1_64 ( .A(asr2_rom_10__0_), .Y(_236_) );
INVX1 INVX1_65 ( .A(asr2_rom_9__0_), .Y(_237_) );
NOR2X1 NOR2X1_31 ( .A(counterdown_counter_2_), .B(_228_), .Y(_238_) );
NAND2X1 NAND2X1_29 ( .A(_238_), .B(_231_), .Y(_239_) );
NAND2X1 NAND2X1_30 ( .A(_233_), .B(_238_), .Y(_240_) );
OAI22X1 OAI22X1_26 ( .A(_236_), .B(_240_), .C(_237_), .D(_239_), .Y(_241_) );
NOR2X1 NOR2X1_32 ( .A(_241_), .B(_235_), .Y(_242_) );
INVX1 INVX1_66 ( .A(asr2_rom_2__0_), .Y(_243_) );
INVX1 INVX1_67 ( .A(asr2_rom_1__0_), .Y(_244_) );
NOR2X1 NOR2X1_33 ( .A(counterdown_counter_3_), .B(counterdown_counter_2_), .Y(_245_) );
NAND2X1 NAND2X1_31 ( .A(_245_), .B(_231_), .Y(_246_) );
NAND2X1 NAND2X1_32 ( .A(_245_), .B(_233_), .Y(_247_) );
OAI22X1 OAI22X1_27 ( .A(_243_), .B(_247_), .C(_244_), .D(_246_), .Y(_248_) );
INVX1 INVX1_68 ( .A(asr2_rom_14__0_), .Y(_249_) );
NAND2X1 NAND2X1_33 ( .A(counterdown_counter_0_), .B(_230_), .Y(_250_) );
NAND2X1 NAND2X1_34 ( .A(counterdown_counter_3_), .B(counterdown_counter_2_), .Y(_251_) );
NOR2X1 NOR2X1_34 ( .A(_251_), .B(_250_), .Y(_252_) );
NAND2X1 NAND2X1_35 ( .A(asr2_rom_13__0_), .B(_252_), .Y(_253_) );
AND2X2 AND2X2_16 ( .A(counterdown_counter_3_), .B(counterdown_counter_2_), .Y(_254_) );
NAND2X1 NAND2X1_36 ( .A(_254_), .B(_233_), .Y(_255_) );
OAI21X1 OAI21X1_9 ( .A(_249_), .B(_255_), .C(_253_), .Y(_256_) );
NOR2X1 NOR2X1_35 ( .A(_248_), .B(_256_), .Y(_257_) );
AND2X2 AND2X2_17 ( .A(counterdown_counter_1_), .B(counterdown_counter_0_), .Y(_258_) );
AND2X2 AND2X2_18 ( .A(_258__bF_buf3), .B(_245_), .Y(_259_) );
NAND2X1 NAND2X1_37 ( .A(asr2_rom_3__0_), .B(_259_), .Y(_260_) );
NOR2X1 NOR2X1_36 ( .A(counterdown_counter_1_), .B(counterdown_counter_0_), .Y(_261_) );
NAND3X1 NAND3X1_65 ( .A(asr2_rom_4__0_), .B(_261__bF_buf3), .C(_229__bF_buf1), .Y(_262_) );
NAND3X1 NAND3X1_66 ( .A(asr2_rom_0__0_), .B(_245_), .C(_261__bF_buf2), .Y(_263_) );
NAND3X1 NAND3X1_67 ( .A(asr2_en_0_), .B(_254_), .C(_258__bF_buf2), .Y(_264_) );
AND2X2 AND2X2_19 ( .A(_264_), .B(_263_), .Y(_265_) );
NAND3X1 NAND3X1_68 ( .A(_260_), .B(_262_), .C(_265_), .Y(_266_) );
NAND3X1 NAND3X1_69 ( .A(asr2_rom_7__0_), .B(_258__bF_buf1), .C(_229__bF_buf0), .Y(_267_) );
NAND3X1 NAND3X1_70 ( .A(asr2_rom_8__0_), .B(_261__bF_buf1), .C(_238_), .Y(_268_) );
NAND2X1 NAND2X1_38 ( .A(counterdown_counter_1_), .B(counterdown_counter_0_), .Y(_269_) );
NOR3X1 NOR3X1_3 ( .A(counterdown_counter_2_), .B(_228_), .C(_269_), .Y(_270_) );
NOR3X1 NOR3X1_4 ( .A(counterdown_counter_1_), .B(counterdown_counter_0_), .C(_251_), .Y(_271_) );
AOI22X1 AOI22X1_9 ( .A(_271_), .B(asr2_rom_12__0_), .C(asr2_rom_11__0_), .D(_270_), .Y(_272_) );
NAND3X1 NAND3X1_71 ( .A(_267_), .B(_268_), .C(_272_), .Y(_273_) );
NOR2X1 NOR2X1_37 ( .A(_266_), .B(_273_), .Y(_274_) );
NAND3X1 NAND3X1_72 ( .A(_242_), .B(_257_), .C(_274_), .Y(asr2_dataout_0_) );
INVX1 INVX1_69 ( .A(asr2_rom_6__1_), .Y(_275_) );
INVX1 INVX1_70 ( .A(asr2_rom_5__1_), .Y(_276_) );
OAI22X1 OAI22X1_28 ( .A(_275_), .B(_234_), .C(_276_), .D(_232_), .Y(_277_) );
INVX1 INVX1_71 ( .A(asr2_rom_10__1_), .Y(_278_) );
INVX1 INVX1_72 ( .A(asr2_rom_9__1_), .Y(_279_) );
OAI22X1 OAI22X1_29 ( .A(_278_), .B(_240_), .C(_279_), .D(_239_), .Y(_280_) );
NOR2X1 NOR2X1_38 ( .A(_280_), .B(_277_), .Y(_281_) );
INVX1 INVX1_73 ( .A(asr2_rom_2__1_), .Y(_282_) );
INVX1 INVX1_74 ( .A(asr2_rom_1__1_), .Y(_283_) );
OAI22X1 OAI22X1_30 ( .A(_282_), .B(_247_), .C(_283_), .D(_246_), .Y(_284_) );
INVX1 INVX1_75 ( .A(asr2_rom_14__1_), .Y(_285_) );
NAND2X1 NAND2X1_39 ( .A(asr2_rom_13__1_), .B(_252_), .Y(_286_) );
OAI21X1 OAI21X1_10 ( .A(_285_), .B(_255_), .C(_286_), .Y(_287_) );
NOR2X1 NOR2X1_39 ( .A(_284_), .B(_287_), .Y(_288_) );
NAND2X1 NAND2X1_40 ( .A(asr2_rom_3__1_), .B(_259_), .Y(_289_) );
NAND3X1 NAND3X1_73 ( .A(asr2_rom_4__1_), .B(_261__bF_buf0), .C(_229__bF_buf3), .Y(_290_) );
NAND3X1 NAND3X1_74 ( .A(asr2_rom_0__1_), .B(_245_), .C(_261__bF_buf3), .Y(_291_) );
NAND3X1 NAND3X1_75 ( .A(asr2_en_1_), .B(_254_), .C(_258__bF_buf0), .Y(_292_) );
AND2X2 AND2X2_20 ( .A(_292_), .B(_291_), .Y(_293_) );
NAND3X1 NAND3X1_76 ( .A(_289_), .B(_290_), .C(_293_), .Y(_294_) );
NAND3X1 NAND3X1_77 ( .A(asr2_rom_7__1_), .B(_258__bF_buf3), .C(_229__bF_buf2), .Y(_295_) );
NAND3X1 NAND3X1_78 ( .A(asr2_rom_8__1_), .B(_261__bF_buf2), .C(_238_), .Y(_296_) );
AOI22X1 AOI22X1_10 ( .A(_271_), .B(asr2_rom_12__1_), .C(asr2_rom_11__1_), .D(_270_), .Y(_297_) );
NAND3X1 NAND3X1_79 ( .A(_295_), .B(_296_), .C(_297_), .Y(_298_) );
NOR2X1 NOR2X1_40 ( .A(_294_), .B(_298_), .Y(_299_) );
NAND3X1 NAND3X1_80 ( .A(_281_), .B(_288_), .C(_299_), .Y(asr2_dataout_1_) );
INVX1 INVX1_76 ( .A(asr2_rom_6__2_), .Y(_300_) );
INVX1 INVX1_77 ( .A(asr2_rom_5__2_), .Y(_301_) );
OAI22X1 OAI22X1_31 ( .A(_300_), .B(_234_), .C(_301_), .D(_232_), .Y(_302_) );
INVX1 INVX1_78 ( .A(asr2_rom_10__2_), .Y(_303_) );
INVX1 INVX1_79 ( .A(asr2_rom_9__2_), .Y(_304_) );
OAI22X1 OAI22X1_32 ( .A(_303_), .B(_240_), .C(_304_), .D(_239_), .Y(_305_) );
NOR2X1 NOR2X1_41 ( .A(_305_), .B(_302_), .Y(_306_) );
INVX1 INVX1_80 ( .A(asr2_rom_2__2_), .Y(_307_) );
INVX1 INVX1_81 ( .A(asr2_rom_1__2_), .Y(_308_) );
OAI22X1 OAI22X1_33 ( .A(_307_), .B(_247_), .C(_308_), .D(_246_), .Y(_309_) );
INVX1 INVX1_82 ( .A(asr2_rom_14__2_), .Y(_310_) );
NAND2X1 NAND2X1_41 ( .A(asr2_rom_13__2_), .B(_252_), .Y(_311_) );
OAI21X1 OAI21X1_11 ( .A(_310_), .B(_255_), .C(_311_), .Y(_312_) );
NOR2X1 NOR2X1_42 ( .A(_309_), .B(_312_), .Y(_313_) );
NAND2X1 NAND2X1_42 ( .A(asr2_rom_3__2_), .B(_259_), .Y(_314_) );
NAND3X1 NAND3X1_81 ( .A(asr2_rom_4__2_), .B(_261__bF_buf1), .C(_229__bF_buf1), .Y(_315_) );
NAND3X1 NAND3X1_82 ( .A(asr2_rom_0__2_), .B(_245_), .C(_261__bF_buf0), .Y(_316_) );
NAND3X1 NAND3X1_83 ( .A(asr2_en_2_), .B(_254_), .C(_258__bF_buf2), .Y(_317_) );
AND2X2 AND2X2_21 ( .A(_317_), .B(_316_), .Y(_318_) );
NAND3X1 NAND3X1_84 ( .A(_314_), .B(_315_), .C(_318_), .Y(_319_) );
NAND3X1 NAND3X1_85 ( .A(asr2_rom_7__2_), .B(_258__bF_buf1), .C(_229__bF_buf0), .Y(_320_) );
NAND3X1 NAND3X1_86 ( .A(asr2_rom_8__2_), .B(_261__bF_buf3), .C(_238_), .Y(_321_) );
AOI22X1 AOI22X1_11 ( .A(_271_), .B(asr2_rom_12__2_), .C(asr2_rom_11__2_), .D(_270_), .Y(_322_) );
NAND3X1 NAND3X1_87 ( .A(_320_), .B(_321_), .C(_322_), .Y(_323_) );
NOR2X1 NOR2X1_43 ( .A(_319_), .B(_323_), .Y(_324_) );
NAND3X1 NAND3X1_88 ( .A(_306_), .B(_313_), .C(_324_), .Y(asr2_dataout_2_) );
INVX1 INVX1_83 ( .A(asr2_rom_6__3_), .Y(_325_) );
INVX1 INVX1_84 ( .A(asr2_rom_5__3_), .Y(_326_) );
OAI22X1 OAI22X1_34 ( .A(_325_), .B(_234_), .C(_326_), .D(_232_), .Y(_327_) );
INVX1 INVX1_85 ( .A(asr2_rom_10__3_), .Y(_328_) );
INVX1 INVX1_86 ( .A(asr2_rom_9__3_), .Y(_329_) );
OAI22X1 OAI22X1_35 ( .A(_328_), .B(_240_), .C(_329_), .D(_239_), .Y(_330_) );
NOR2X1 NOR2X1_44 ( .A(_330_), .B(_327_), .Y(_331_) );
INVX1 INVX1_87 ( .A(asr2_rom_2__3_), .Y(_332_) );
INVX1 INVX1_88 ( .A(asr2_rom_1__3_), .Y(_333_) );
OAI22X1 OAI22X1_36 ( .A(_332_), .B(_247_), .C(_333_), .D(_246_), .Y(_334_) );
INVX1 INVX1_89 ( .A(asr2_rom_14__3_), .Y(_335_) );
NAND2X1 NAND2X1_43 ( .A(asr2_rom_13__3_), .B(_252_), .Y(_336_) );
OAI21X1 OAI21X1_12 ( .A(_335_), .B(_255_), .C(_336_), .Y(_337_) );
NOR2X1 NOR2X1_45 ( .A(_334_), .B(_337_), .Y(_338_) );
NAND2X1 NAND2X1_44 ( .A(asr2_rom_3__3_), .B(_259_), .Y(_339_) );
NAND3X1 NAND3X1_89 ( .A(asr2_rom_4__3_), .B(_261__bF_buf2), .C(_229__bF_buf3), .Y(_340_) );
NAND3X1 NAND3X1_90 ( .A(asr2_rom_0__3_), .B(_245_), .C(_261__bF_buf1), .Y(_341_) );
NAND3X1 NAND3X1_91 ( .A(asr2_en_3_), .B(_254_), .C(_258__bF_buf0), .Y(_342_) );
AND2X2 AND2X2_22 ( .A(_342_), .B(_341_), .Y(_343_) );
NAND3X1 NAND3X1_92 ( .A(_339_), .B(_340_), .C(_343_), .Y(_344_) );
NAND3X1 NAND3X1_93 ( .A(asr2_rom_7__3_), .B(_258__bF_buf3), .C(_229__bF_buf2), .Y(_345_) );
NAND3X1 NAND3X1_94 ( .A(asr2_rom_8__3_), .B(_261__bF_buf0), .C(_238_), .Y(_346_) );
AOI22X1 AOI22X1_12 ( .A(_271_), .B(asr2_rom_12__3_), .C(asr2_rom_11__3_), .D(_270_), .Y(_347_) );
NAND3X1 NAND3X1_95 ( .A(_345_), .B(_346_), .C(_347_), .Y(_348_) );
NOR2X1 NOR2X1_46 ( .A(_344_), .B(_348_), .Y(_349_) );
NAND3X1 NAND3X1_96 ( .A(_331_), .B(_338_), .C(_349_), .Y(asr2_dataout_3_) );
INVX1 INVX1_90 ( .A(asr2_rom_6__4_), .Y(_350_) );
INVX1 INVX1_91 ( .A(asr2_rom_5__4_), .Y(_351_) );
OAI22X1 OAI22X1_37 ( .A(_350_), .B(_234_), .C(_351_), .D(_232_), .Y(_352_) );
INVX1 INVX1_92 ( .A(asr2_rom_10__4_), .Y(_353_) );
INVX1 INVX1_93 ( .A(asr2_rom_9__4_), .Y(_354_) );
OAI22X1 OAI22X1_38 ( .A(_353_), .B(_240_), .C(_354_), .D(_239_), .Y(_355_) );
NOR2X1 NOR2X1_47 ( .A(_355_), .B(_352_), .Y(_356_) );
INVX1 INVX1_94 ( .A(asr2_rom_2__4_), .Y(_357_) );
INVX1 INVX1_95 ( .A(asr2_rom_1__4_), .Y(_358_) );
OAI22X1 OAI22X1_39 ( .A(_357_), .B(_247_), .C(_358_), .D(_246_), .Y(_359_) );
INVX1 INVX1_96 ( .A(asr2_rom_14__4_), .Y(_360_) );
NAND2X1 NAND2X1_45 ( .A(asr2_rom_13__4_), .B(_252_), .Y(_361_) );
OAI21X1 OAI21X1_13 ( .A(_360_), .B(_255_), .C(_361_), .Y(_362_) );
NOR2X1 NOR2X1_48 ( .A(_359_), .B(_362_), .Y(_363_) );
NAND2X1 NAND2X1_46 ( .A(asr2_rom_3__4_), .B(_259_), .Y(_364_) );
NAND3X1 NAND3X1_97 ( .A(asr2_rom_4__4_), .B(_261__bF_buf3), .C(_229__bF_buf1), .Y(_365_) );
NAND3X1 NAND3X1_98 ( .A(asr2_rom_0__4_), .B(_245_), .C(_261__bF_buf2), .Y(_366_) );
NAND3X1 NAND3X1_99 ( .A(asr2_en_4_), .B(_254_), .C(_258__bF_buf2), .Y(_367_) );
AND2X2 AND2X2_23 ( .A(_367_), .B(_366_), .Y(_368_) );
NAND3X1 NAND3X1_100 ( .A(_364_), .B(_365_), .C(_368_), .Y(_369_) );
NAND3X1 NAND3X1_101 ( .A(asr2_rom_7__4_), .B(_258__bF_buf1), .C(_229__bF_buf0), .Y(_370_) );
NAND3X1 NAND3X1_102 ( .A(asr2_rom_8__4_), .B(_261__bF_buf1), .C(_238_), .Y(_371_) );
AOI22X1 AOI22X1_13 ( .A(_271_), .B(asr2_rom_12__4_), .C(asr2_rom_11__4_), .D(_270_), .Y(_372_) );
NAND3X1 NAND3X1_103 ( .A(_370_), .B(_371_), .C(_372_), .Y(_373_) );
NOR2X1 NOR2X1_49 ( .A(_369_), .B(_373_), .Y(_374_) );
NAND3X1 NAND3X1_104 ( .A(_356_), .B(_363_), .C(_374_), .Y(asr2_dataout_4_) );
INVX1 INVX1_97 ( .A(asr2_rom_6__5_), .Y(_375_) );
INVX1 INVX1_98 ( .A(asr2_rom_5__5_), .Y(_376_) );
OAI22X1 OAI22X1_40 ( .A(_375_), .B(_234_), .C(_376_), .D(_232_), .Y(_377_) );
INVX1 INVX1_99 ( .A(asr2_rom_10__5_), .Y(_378_) );
INVX1 INVX1_100 ( .A(asr2_rom_9__5_), .Y(_379_) );
OAI22X1 OAI22X1_41 ( .A(_378_), .B(_240_), .C(_379_), .D(_239_), .Y(_380_) );
NOR2X1 NOR2X1_50 ( .A(_380_), .B(_377_), .Y(_381_) );
INVX1 INVX1_101 ( .A(asr2_rom_2__5_), .Y(_382_) );
INVX1 INVX1_102 ( .A(asr2_rom_1__5_), .Y(_383_) );
OAI22X1 OAI22X1_42 ( .A(_382_), .B(_247_), .C(_383_), .D(_246_), .Y(_384_) );
INVX1 INVX1_103 ( .A(asr2_rom_14__5_), .Y(_385_) );
NAND2X1 NAND2X1_47 ( .A(asr2_rom_13__5_), .B(_252_), .Y(_386_) );
OAI21X1 OAI21X1_14 ( .A(_385_), .B(_255_), .C(_386_), .Y(_387_) );
NOR2X1 NOR2X1_51 ( .A(_384_), .B(_387_), .Y(_388_) );
NAND2X1 NAND2X1_48 ( .A(asr2_rom_3__5_), .B(_259_), .Y(_389_) );
NAND3X1 NAND3X1_105 ( .A(asr2_rom_4__5_), .B(_261__bF_buf0), .C(_229__bF_buf3), .Y(_390_) );
NAND3X1 NAND3X1_106 ( .A(asr2_rom_0__5_), .B(_245_), .C(_261__bF_buf3), .Y(_391_) );
NAND3X1 NAND3X1_107 ( .A(asr2_en_5_), .B(_254_), .C(_258__bF_buf0), .Y(_392_) );
AND2X2 AND2X2_24 ( .A(_392_), .B(_391_), .Y(_393_) );
NAND3X1 NAND3X1_108 ( .A(_389_), .B(_390_), .C(_393_), .Y(_394_) );
NAND3X1 NAND3X1_109 ( .A(asr2_rom_7__5_), .B(_258__bF_buf3), .C(_229__bF_buf2), .Y(_395_) );
NAND3X1 NAND3X1_110 ( .A(asr2_rom_8__5_), .B(_261__bF_buf2), .C(_238_), .Y(_396_) );
AOI22X1 AOI22X1_14 ( .A(_271_), .B(asr2_rom_12__5_), .C(asr2_rom_11__5_), .D(_270_), .Y(_397_) );
NAND3X1 NAND3X1_111 ( .A(_395_), .B(_396_), .C(_397_), .Y(_398_) );
NOR2X1 NOR2X1_52 ( .A(_394_), .B(_398_), .Y(_399_) );
NAND3X1 NAND3X1_112 ( .A(_381_), .B(_388_), .C(_399_), .Y(asr2_dataout_5_) );
INVX1 INVX1_104 ( .A(asr2_rom_6__6_), .Y(_400_) );
INVX1 INVX1_105 ( .A(asr2_rom_5__6_), .Y(_401_) );
OAI22X1 OAI22X1_43 ( .A(_400_), .B(_234_), .C(_401_), .D(_232_), .Y(_402_) );
INVX1 INVX1_106 ( .A(asr2_rom_10__6_), .Y(_403_) );
INVX1 INVX1_107 ( .A(asr2_rom_9__6_), .Y(_404_) );
OAI22X1 OAI22X1_44 ( .A(_403_), .B(_240_), .C(_404_), .D(_239_), .Y(_405_) );
NOR2X1 NOR2X1_53 ( .A(_405_), .B(_402_), .Y(_406_) );
INVX1 INVX1_108 ( .A(asr2_rom_2__6_), .Y(_407_) );
INVX1 INVX1_109 ( .A(asr2_rom_1__6_), .Y(_408_) );
OAI22X1 OAI22X1_45 ( .A(_407_), .B(_247_), .C(_408_), .D(_246_), .Y(_409_) );
INVX1 INVX1_110 ( .A(asr2_rom_14__6_), .Y(_410_) );
NAND2X1 NAND2X1_49 ( .A(asr2_rom_13__6_), .B(_252_), .Y(_411_) );
OAI21X1 OAI21X1_15 ( .A(_410_), .B(_255_), .C(_411_), .Y(_412_) );
NOR2X1 NOR2X1_54 ( .A(_409_), .B(_412_), .Y(_413_) );
NAND2X1 NAND2X1_50 ( .A(asr2_rom_3__6_), .B(_259_), .Y(_414_) );
NAND3X1 NAND3X1_113 ( .A(asr2_rom_4__6_), .B(_261__bF_buf1), .C(_229__bF_buf1), .Y(_415_) );
NAND3X1 NAND3X1_114 ( .A(asr2_rom_0__6_), .B(_245_), .C(_261__bF_buf0), .Y(_416_) );
NAND3X1 NAND3X1_115 ( .A(asr2_en_6_), .B(_254_), .C(_258__bF_buf2), .Y(_417_) );
AND2X2 AND2X2_25 ( .A(_417_), .B(_416_), .Y(_418_) );
NAND3X1 NAND3X1_116 ( .A(_414_), .B(_415_), .C(_418_), .Y(_419_) );
NAND3X1 NAND3X1_117 ( .A(asr2_rom_7__6_), .B(_258__bF_buf1), .C(_229__bF_buf0), .Y(_420_) );
NAND3X1 NAND3X1_118 ( .A(asr2_rom_8__6_), .B(_261__bF_buf3), .C(_238_), .Y(_421_) );
AOI22X1 AOI22X1_15 ( .A(_271_), .B(asr2_rom_12__6_), .C(asr2_rom_11__6_), .D(_270_), .Y(_422_) );
NAND3X1 NAND3X1_119 ( .A(_420_), .B(_421_), .C(_422_), .Y(_423_) );
NOR2X1 NOR2X1_55 ( .A(_419_), .B(_423_), .Y(_424_) );
NAND3X1 NAND3X1_120 ( .A(_406_), .B(_413_), .C(_424_), .Y(asr2_dataout_6_) );
INVX1 INVX1_111 ( .A(asr2_rom_6__7_), .Y(_425_) );
INVX1 INVX1_112 ( .A(asr2_rom_5__7_), .Y(_426_) );
OAI22X1 OAI22X1_46 ( .A(_425_), .B(_234_), .C(_426_), .D(_232_), .Y(_427_) );
INVX1 INVX1_113 ( .A(asr2_rom_10__7_), .Y(_428_) );
INVX1 INVX1_114 ( .A(asr2_rom_9__7_), .Y(_429_) );
OAI22X1 OAI22X1_47 ( .A(_428_), .B(_240_), .C(_429_), .D(_239_), .Y(_430_) );
NOR2X1 NOR2X1_56 ( .A(_430_), .B(_427_), .Y(_431_) );
INVX1 INVX1_115 ( .A(asr2_rom_2__7_), .Y(_432_) );
INVX1 INVX1_116 ( .A(asr2_rom_1__7_), .Y(_433_) );
OAI22X1 OAI22X1_48 ( .A(_432_), .B(_247_), .C(_433_), .D(_246_), .Y(_434_) );
INVX1 INVX1_117 ( .A(asr2_rom_14__7_), .Y(_435_) );
NAND2X1 NAND2X1_51 ( .A(asr2_rom_13__7_), .B(_252_), .Y(_436_) );
OAI21X1 OAI21X1_16 ( .A(_435_), .B(_255_), .C(_436_), .Y(_437_) );
NOR2X1 NOR2X1_57 ( .A(_434_), .B(_437_), .Y(_438_) );
NAND2X1 NAND2X1_52 ( .A(asr2_rom_3__7_), .B(_259_), .Y(_439_) );
NAND3X1 NAND3X1_121 ( .A(asr2_rom_4__7_), .B(_261__bF_buf2), .C(_229__bF_buf3), .Y(_440_) );
NAND3X1 NAND3X1_122 ( .A(asr2_rom_0__7_), .B(_245_), .C(_261__bF_buf1), .Y(_441_) );
NAND3X1 NAND3X1_123 ( .A(asr2_en_7_), .B(_254_), .C(_258__bF_buf0), .Y(_442_) );
AND2X2 AND2X2_26 ( .A(_442_), .B(_441_), .Y(_443_) );
NAND3X1 NAND3X1_124 ( .A(_439_), .B(_440_), .C(_443_), .Y(_444_) );
NAND3X1 NAND3X1_125 ( .A(asr2_rom_7__7_), .B(_258__bF_buf3), .C(_229__bF_buf2), .Y(_445_) );
NAND3X1 NAND3X1_126 ( .A(asr2_rom_8__7_), .B(_261__bF_buf0), .C(_238_), .Y(_446_) );
AOI22X1 AOI22X1_16 ( .A(_271_), .B(asr2_rom_12__7_), .C(asr2_rom_11__7_), .D(_270_), .Y(_447_) );
NAND3X1 NAND3X1_127 ( .A(_445_), .B(_446_), .C(_447_), .Y(_448_) );
NOR2X1 NOR2X1_58 ( .A(_444_), .B(_448_), .Y(_449_) );
NAND3X1 NAND3X1_128 ( .A(_431_), .B(_438_), .C(_449_), .Y(asr2_dataout_7_) );
INVX1 INVX1_118 ( .A(rst_bF_buf4), .Y(_225_) );
DFFSR DFFSR_129 ( .CLK(clk2_clkout_bF_buf39), .D(asr1_en_0_), .Q(asr2_rom_0__0_), .R(_225__bF_buf10), .S(vdd) );
DFFSR DFFSR_130 ( .CLK(clk2_clkout_bF_buf38), .D(asr1_en_1_), .Q(asr2_rom_0__1_), .R(_225__bF_buf9), .S(vdd) );
DFFSR DFFSR_131 ( .CLK(clk2_clkout_bF_buf37), .D(asr1_en_2_), .Q(asr2_rom_0__2_), .R(_225__bF_buf8), .S(vdd) );
DFFSR DFFSR_132 ( .CLK(clk2_clkout_bF_buf36), .D(asr1_en_3_), .Q(asr2_rom_0__3_), .R(_225__bF_buf7), .S(vdd) );
DFFSR DFFSR_133 ( .CLK(clk2_clkout_bF_buf35), .D(asr1_en_4_), .Q(asr2_rom_0__4_), .R(_225__bF_buf6), .S(vdd) );
DFFSR DFFSR_134 ( .CLK(clk2_clkout_bF_buf34), .D(asr1_en_5_), .Q(asr2_rom_0__5_), .R(_225__bF_buf5), .S(vdd) );
DFFSR DFFSR_135 ( .CLK(clk2_clkout_bF_buf33), .D(asr1_en_6_), .Q(asr2_rom_0__6_), .R(_225__bF_buf4), .S(vdd) );
DFFSR DFFSR_136 ( .CLK(clk2_clkout_bF_buf32), .D(asr1_en_7_), .Q(asr2_rom_0__7_), .R(_225__bF_buf3), .S(vdd) );
DFFSR DFFSR_137 ( .CLK(clk2_clkout_bF_buf31), .D(asr2_rom_6__0_), .Q(asr2_rom_7__0_), .R(_225__bF_buf2), .S(vdd) );
DFFSR DFFSR_138 ( .CLK(clk2_clkout_bF_buf30), .D(asr2_rom_6__1_), .Q(asr2_rom_7__1_), .R(_225__bF_buf1), .S(vdd) );
DFFSR DFFSR_139 ( .CLK(clk2_clkout_bF_buf29), .D(asr2_rom_6__2_), .Q(asr2_rom_7__2_), .R(_225__bF_buf0), .S(vdd) );
DFFSR DFFSR_140 ( .CLK(clk2_clkout_bF_buf28), .D(asr2_rom_6__3_), .Q(asr2_rom_7__3_), .R(_225__bF_buf10), .S(vdd) );
DFFSR DFFSR_141 ( .CLK(clk2_clkout_bF_buf27), .D(asr2_rom_6__4_), .Q(asr2_rom_7__4_), .R(_225__bF_buf9), .S(vdd) );
DFFSR DFFSR_142 ( .CLK(clk2_clkout_bF_buf26), .D(asr2_rom_6__5_), .Q(asr2_rom_7__5_), .R(_225__bF_buf8), .S(vdd) );
DFFSR DFFSR_143 ( .CLK(clk2_clkout_bF_buf25), .D(asr2_rom_6__6_), .Q(asr2_rom_7__6_), .R(_225__bF_buf7), .S(vdd) );
DFFSR DFFSR_144 ( .CLK(clk2_clkout_bF_buf24), .D(asr2_rom_6__7_), .Q(asr2_rom_7__7_), .R(_225__bF_buf6), .S(vdd) );
DFFSR DFFSR_145 ( .CLK(clk2_clkout_bF_buf23), .D(asr2_rom_1__0_), .Q(asr2_rom_2__0_), .R(_225__bF_buf5), .S(vdd) );
DFFSR DFFSR_146 ( .CLK(clk2_clkout_bF_buf22), .D(asr2_rom_1__1_), .Q(asr2_rom_2__1_), .R(_225__bF_buf4), .S(vdd) );
DFFSR DFFSR_147 ( .CLK(clk2_clkout_bF_buf21), .D(asr2_rom_1__2_), .Q(asr2_rom_2__2_), .R(_225__bF_buf3), .S(vdd) );
DFFSR DFFSR_148 ( .CLK(clk2_clkout_bF_buf20), .D(asr2_rom_1__3_), .Q(asr2_rom_2__3_), .R(_225__bF_buf2), .S(vdd) );
DFFSR DFFSR_149 ( .CLK(clk2_clkout_bF_buf19), .D(asr2_rom_1__4_), .Q(asr2_rom_2__4_), .R(_225__bF_buf1), .S(vdd) );
DFFSR DFFSR_150 ( .CLK(clk2_clkout_bF_buf18), .D(asr2_rom_1__5_), .Q(asr2_rom_2__5_), .R(_225__bF_buf0), .S(vdd) );
DFFSR DFFSR_151 ( .CLK(clk2_clkout_bF_buf17), .D(asr2_rom_1__6_), .Q(asr2_rom_2__6_), .R(_225__bF_buf10), .S(vdd) );
DFFSR DFFSR_152 ( .CLK(clk2_clkout_bF_buf16), .D(asr2_rom_1__7_), .Q(asr2_rom_2__7_), .R(_225__bF_buf9), .S(vdd) );
DFFSR DFFSR_153 ( .CLK(clk2_clkout_bF_buf15), .D(asr2_rom_0__0_), .Q(asr2_rom_1__0_), .R(_225__bF_buf8), .S(vdd) );
DFFSR DFFSR_154 ( .CLK(clk2_clkout_bF_buf14), .D(asr2_rom_0__1_), .Q(asr2_rom_1__1_), .R(_225__bF_buf7), .S(vdd) );
DFFSR DFFSR_155 ( .CLK(clk2_clkout_bF_buf13), .D(asr2_rom_0__2_), .Q(asr2_rom_1__2_), .R(_225__bF_buf6), .S(vdd) );
DFFSR DFFSR_156 ( .CLK(clk2_clkout_bF_buf12), .D(asr2_rom_0__3_), .Q(asr2_rom_1__3_), .R(_225__bF_buf5), .S(vdd) );
DFFSR DFFSR_157 ( .CLK(clk2_clkout_bF_buf11), .D(asr2_rom_0__4_), .Q(asr2_rom_1__4_), .R(_225__bF_buf4), .S(vdd) );
DFFSR DFFSR_158 ( .CLK(clk2_clkout_bF_buf10), .D(asr2_rom_0__5_), .Q(asr2_rom_1__5_), .R(_225__bF_buf3), .S(vdd) );
DFFSR DFFSR_159 ( .CLK(clk2_clkout_bF_buf9), .D(asr2_rom_0__6_), .Q(asr2_rom_1__6_), .R(_225__bF_buf2), .S(vdd) );
DFFSR DFFSR_160 ( .CLK(clk2_clkout_bF_buf8), .D(asr2_rom_0__7_), .Q(asr2_rom_1__7_), .R(_225__bF_buf1), .S(vdd) );
DFFSR DFFSR_161 ( .CLK(clk2_clkout_bF_buf7), .D(asr2_rom_2__0_), .Q(asr2_rom_3__0_), .R(_225__bF_buf0), .S(vdd) );
DFFSR DFFSR_162 ( .CLK(clk2_clkout_bF_buf6), .D(asr2_rom_2__1_), .Q(asr2_rom_3__1_), .R(_225__bF_buf10), .S(vdd) );
DFFSR DFFSR_163 ( .CLK(clk2_clkout_bF_buf5), .D(asr2_rom_2__2_), .Q(asr2_rom_3__2_), .R(_225__bF_buf9), .S(vdd) );
DFFSR DFFSR_164 ( .CLK(clk2_clkout_bF_buf4), .D(asr2_rom_2__3_), .Q(asr2_rom_3__3_), .R(_225__bF_buf8), .S(vdd) );
DFFSR DFFSR_165 ( .CLK(clk2_clkout_bF_buf3), .D(asr2_rom_2__4_), .Q(asr2_rom_3__4_), .R(_225__bF_buf7), .S(vdd) );
DFFSR DFFSR_166 ( .CLK(clk2_clkout_bF_buf2), .D(asr2_rom_2__5_), .Q(asr2_rom_3__5_), .R(_225__bF_buf6), .S(vdd) );
DFFSR DFFSR_167 ( .CLK(clk2_clkout_bF_buf1), .D(asr2_rom_2__6_), .Q(asr2_rom_3__6_), .R(_225__bF_buf5), .S(vdd) );
DFFSR DFFSR_168 ( .CLK(clk2_clkout_bF_buf0), .D(asr2_rom_2__7_), .Q(asr2_rom_3__7_), .R(_225__bF_buf4), .S(vdd) );
DFFSR DFFSR_169 ( .CLK(clk2_clkout_bF_buf41), .D(asr2_rom_3__0_), .Q(asr2_rom_4__0_), .R(_225__bF_buf3), .S(vdd) );
DFFSR DFFSR_170 ( .CLK(clk2_clkout_bF_buf40), .D(asr2_rom_3__1_), .Q(asr2_rom_4__1_), .R(_225__bF_buf2), .S(vdd) );
DFFSR DFFSR_171 ( .CLK(clk2_clkout_bF_buf39), .D(asr2_rom_3__2_), .Q(asr2_rom_4__2_), .R(_225__bF_buf1), .S(vdd) );
DFFSR DFFSR_172 ( .CLK(clk2_clkout_bF_buf38), .D(asr2_rom_3__3_), .Q(asr2_rom_4__3_), .R(_225__bF_buf0), .S(vdd) );
DFFSR DFFSR_173 ( .CLK(clk2_clkout_bF_buf37), .D(asr2_rom_3__4_), .Q(asr2_rom_4__4_), .R(_225__bF_buf10), .S(vdd) );
DFFSR DFFSR_174 ( .CLK(clk2_clkout_bF_buf36), .D(asr2_rom_3__5_), .Q(asr2_rom_4__5_), .R(_225__bF_buf9), .S(vdd) );
DFFSR DFFSR_175 ( .CLK(clk2_clkout_bF_buf35), .D(asr2_rom_3__6_), .Q(asr2_rom_4__6_), .R(_225__bF_buf8), .S(vdd) );
DFFSR DFFSR_176 ( .CLK(clk2_clkout_bF_buf34), .D(asr2_rom_3__7_), .Q(asr2_rom_4__7_), .R(_225__bF_buf7), .S(vdd) );
DFFSR DFFSR_177 ( .CLK(clk2_clkout_bF_buf33), .D(asr2_rom_5__0_), .Q(asr2_rom_6__0_), .R(_225__bF_buf6), .S(vdd) );
DFFSR DFFSR_178 ( .CLK(clk2_clkout_bF_buf32), .D(asr2_rom_5__1_), .Q(asr2_rom_6__1_), .R(_225__bF_buf5), .S(vdd) );
DFFSR DFFSR_179 ( .CLK(clk2_clkout_bF_buf31), .D(asr2_rom_5__2_), .Q(asr2_rom_6__2_), .R(_225__bF_buf4), .S(vdd) );
DFFSR DFFSR_180 ( .CLK(clk2_clkout_bF_buf30), .D(asr2_rom_5__3_), .Q(asr2_rom_6__3_), .R(_225__bF_buf3), .S(vdd) );
DFFSR DFFSR_181 ( .CLK(clk2_clkout_bF_buf29), .D(asr2_rom_5__4_), .Q(asr2_rom_6__4_), .R(_225__bF_buf2), .S(vdd) );
DFFSR DFFSR_182 ( .CLK(clk2_clkout_bF_buf28), .D(asr2_rom_5__5_), .Q(asr2_rom_6__5_), .R(_225__bF_buf1), .S(vdd) );
DFFSR DFFSR_183 ( .CLK(clk2_clkout_bF_buf27), .D(asr2_rom_5__6_), .Q(asr2_rom_6__6_), .R(_225__bF_buf0), .S(vdd) );
DFFSR DFFSR_184 ( .CLK(clk2_clkout_bF_buf26), .D(asr2_rom_5__7_), .Q(asr2_rom_6__7_), .R(_225__bF_buf10), .S(vdd) );
DFFSR DFFSR_185 ( .CLK(clk2_clkout_bF_buf25), .D(asr2_rom_4__0_), .Q(asr2_rom_5__0_), .R(_225__bF_buf9), .S(vdd) );
DFFSR DFFSR_186 ( .CLK(clk2_clkout_bF_buf24), .D(asr2_rom_4__1_), .Q(asr2_rom_5__1_), .R(_225__bF_buf8), .S(vdd) );
DFFSR DFFSR_187 ( .CLK(clk2_clkout_bF_buf23), .D(asr2_rom_4__2_), .Q(asr2_rom_5__2_), .R(_225__bF_buf7), .S(vdd) );
DFFSR DFFSR_188 ( .CLK(clk2_clkout_bF_buf22), .D(asr2_rom_4__3_), .Q(asr2_rom_5__3_), .R(_225__bF_buf6), .S(vdd) );
DFFSR DFFSR_189 ( .CLK(clk2_clkout_bF_buf21), .D(asr2_rom_4__4_), .Q(asr2_rom_5__4_), .R(_225__bF_buf5), .S(vdd) );
DFFSR DFFSR_190 ( .CLK(clk2_clkout_bF_buf20), .D(asr2_rom_4__5_), .Q(asr2_rom_5__5_), .R(_225__bF_buf4), .S(vdd) );
DFFSR DFFSR_191 ( .CLK(clk2_clkout_bF_buf19), .D(asr2_rom_4__6_), .Q(asr2_rom_5__6_), .R(_225__bF_buf3), .S(vdd) );
DFFSR DFFSR_192 ( .CLK(clk2_clkout_bF_buf18), .D(asr2_rom_4__7_), .Q(asr2_rom_5__7_), .R(_225__bF_buf2), .S(vdd) );
DFFSR DFFSR_193 ( .CLK(clk2_clkout_bF_buf17), .D(asr2_rom_7__0_), .Q(asr2_rom_8__0_), .R(_225__bF_buf1), .S(vdd) );
DFFSR DFFSR_194 ( .CLK(clk2_clkout_bF_buf16), .D(asr2_rom_7__1_), .Q(asr2_rom_8__1_), .R(_225__bF_buf0), .S(vdd) );
DFFSR DFFSR_195 ( .CLK(clk2_clkout_bF_buf15), .D(asr2_rom_7__2_), .Q(asr2_rom_8__2_), .R(_225__bF_buf10), .S(vdd) );
DFFSR DFFSR_196 ( .CLK(clk2_clkout_bF_buf14), .D(asr2_rom_7__3_), .Q(asr2_rom_8__3_), .R(_225__bF_buf9), .S(vdd) );
DFFSR DFFSR_197 ( .CLK(clk2_clkout_bF_buf13), .D(asr2_rom_7__4_), .Q(asr2_rom_8__4_), .R(_225__bF_buf8), .S(vdd) );
DFFSR DFFSR_198 ( .CLK(clk2_clkout_bF_buf12), .D(asr2_rom_7__5_), .Q(asr2_rom_8__5_), .R(_225__bF_buf7), .S(vdd) );
DFFSR DFFSR_199 ( .CLK(clk2_clkout_bF_buf11), .D(asr2_rom_7__6_), .Q(asr2_rom_8__6_), .R(_225__bF_buf6), .S(vdd) );
DFFSR DFFSR_200 ( .CLK(clk2_clkout_bF_buf10), .D(asr2_rom_7__7_), .Q(asr2_rom_8__7_), .R(_225__bF_buf5), .S(vdd) );
DFFSR DFFSR_201 ( .CLK(clk2_clkout_bF_buf9), .D(asr2_rom_8__0_), .Q(asr2_rom_9__0_), .R(_225__bF_buf4), .S(vdd) );
DFFSR DFFSR_202 ( .CLK(clk2_clkout_bF_buf8), .D(asr2_rom_8__1_), .Q(asr2_rom_9__1_), .R(_225__bF_buf3), .S(vdd) );
DFFSR DFFSR_203 ( .CLK(clk2_clkout_bF_buf7), .D(asr2_rom_8__2_), .Q(asr2_rom_9__2_), .R(_225__bF_buf2), .S(vdd) );
DFFSR DFFSR_204 ( .CLK(clk2_clkout_bF_buf6), .D(asr2_rom_8__3_), .Q(asr2_rom_9__3_), .R(_225__bF_buf1), .S(vdd) );
DFFSR DFFSR_205 ( .CLK(clk2_clkout_bF_buf5), .D(asr2_rom_8__4_), .Q(asr2_rom_9__4_), .R(_225__bF_buf0), .S(vdd) );
DFFSR DFFSR_206 ( .CLK(clk2_clkout_bF_buf4), .D(asr2_rom_8__5_), .Q(asr2_rom_9__5_), .R(_225__bF_buf10), .S(vdd) );
DFFSR DFFSR_207 ( .CLK(clk2_clkout_bF_buf3), .D(asr2_rom_8__6_), .Q(asr2_rom_9__6_), .R(_225__bF_buf9), .S(vdd) );
DFFSR DFFSR_208 ( .CLK(clk2_clkout_bF_buf2), .D(asr2_rom_8__7_), .Q(asr2_rom_9__7_), .R(_225__bF_buf8), .S(vdd) );
DFFSR DFFSR_209 ( .CLK(clk2_clkout_bF_buf1), .D(asr2_rom_9__0_), .Q(asr2_rom_10__0_), .R(_225__bF_buf7), .S(vdd) );
DFFSR DFFSR_210 ( .CLK(clk2_clkout_bF_buf0), .D(asr2_rom_9__1_), .Q(asr2_rom_10__1_), .R(_225__bF_buf6), .S(vdd) );
DFFSR DFFSR_211 ( .CLK(clk2_clkout_bF_buf41), .D(asr2_rom_9__2_), .Q(asr2_rom_10__2_), .R(_225__bF_buf5), .S(vdd) );
DFFSR DFFSR_212 ( .CLK(clk2_clkout_bF_buf40), .D(asr2_rom_9__3_), .Q(asr2_rom_10__3_), .R(_225__bF_buf4), .S(vdd) );
DFFSR DFFSR_213 ( .CLK(clk2_clkout_bF_buf39), .D(asr2_rom_9__4_), .Q(asr2_rom_10__4_), .R(_225__bF_buf3), .S(vdd) );
DFFSR DFFSR_214 ( .CLK(clk2_clkout_bF_buf38), .D(asr2_rom_9__5_), .Q(asr2_rom_10__5_), .R(_225__bF_buf2), .S(vdd) );
DFFSR DFFSR_215 ( .CLK(clk2_clkout_bF_buf37), .D(asr2_rom_9__6_), .Q(asr2_rom_10__6_), .R(_225__bF_buf1), .S(vdd) );
DFFSR DFFSR_216 ( .CLK(clk2_clkout_bF_buf36), .D(asr2_rom_9__7_), .Q(asr2_rom_10__7_), .R(_225__bF_buf0), .S(vdd) );
DFFSR DFFSR_217 ( .CLK(clk2_clkout_bF_buf35), .D(asr2_rom_10__0_), .Q(asr2_rom_11__0_), .R(_225__bF_buf10), .S(vdd) );
DFFSR DFFSR_218 ( .CLK(clk2_clkout_bF_buf34), .D(asr2_rom_10__1_), .Q(asr2_rom_11__1_), .R(_225__bF_buf9), .S(vdd) );
DFFSR DFFSR_219 ( .CLK(clk2_clkout_bF_buf33), .D(asr2_rom_10__2_), .Q(asr2_rom_11__2_), .R(_225__bF_buf8), .S(vdd) );
DFFSR DFFSR_220 ( .CLK(clk2_clkout_bF_buf32), .D(asr2_rom_10__3_), .Q(asr2_rom_11__3_), .R(_225__bF_buf7), .S(vdd) );
DFFSR DFFSR_221 ( .CLK(clk2_clkout_bF_buf31), .D(asr2_rom_10__4_), .Q(asr2_rom_11__4_), .R(_225__bF_buf6), .S(vdd) );
DFFSR DFFSR_222 ( .CLK(clk2_clkout_bF_buf30), .D(asr2_rom_10__5_), .Q(asr2_rom_11__5_), .R(_225__bF_buf5), .S(vdd) );
DFFSR DFFSR_223 ( .CLK(clk2_clkout_bF_buf29), .D(asr2_rom_10__6_), .Q(asr2_rom_11__6_), .R(_225__bF_buf4), .S(vdd) );
DFFSR DFFSR_224 ( .CLK(clk2_clkout_bF_buf28), .D(asr2_rom_10__7_), .Q(asr2_rom_11__7_), .R(_225__bF_buf3), .S(vdd) );
DFFSR DFFSR_225 ( .CLK(clk2_clkout_bF_buf27), .D(asr2_rom_11__0_), .Q(asr2_rom_12__0_), .R(_225__bF_buf2), .S(vdd) );
DFFSR DFFSR_226 ( .CLK(clk2_clkout_bF_buf26), .D(asr2_rom_11__1_), .Q(asr2_rom_12__1_), .R(_225__bF_buf1), .S(vdd) );
DFFSR DFFSR_227 ( .CLK(clk2_clkout_bF_buf25), .D(asr2_rom_11__2_), .Q(asr2_rom_12__2_), .R(_225__bF_buf0), .S(vdd) );
DFFSR DFFSR_228 ( .CLK(clk2_clkout_bF_buf24), .D(asr2_rom_11__3_), .Q(asr2_rom_12__3_), .R(_225__bF_buf10), .S(vdd) );
DFFSR DFFSR_229 ( .CLK(clk2_clkout_bF_buf23), .D(asr2_rom_11__4_), .Q(asr2_rom_12__4_), .R(_225__bF_buf9), .S(vdd) );
DFFSR DFFSR_230 ( .CLK(clk2_clkout_bF_buf22), .D(asr2_rom_11__5_), .Q(asr2_rom_12__5_), .R(_225__bF_buf8), .S(vdd) );
DFFSR DFFSR_231 ( .CLK(clk2_clkout_bF_buf21), .D(asr2_rom_11__6_), .Q(asr2_rom_12__6_), .R(_225__bF_buf7), .S(vdd) );
DFFSR DFFSR_232 ( .CLK(clk2_clkout_bF_buf20), .D(asr2_rom_11__7_), .Q(asr2_rom_12__7_), .R(_225__bF_buf6), .S(vdd) );
DFFSR DFFSR_233 ( .CLK(clk2_clkout_bF_buf19), .D(asr2_rom_12__0_), .Q(asr2_rom_13__0_), .R(_225__bF_buf5), .S(vdd) );
DFFSR DFFSR_234 ( .CLK(clk2_clkout_bF_buf18), .D(asr2_rom_12__1_), .Q(asr2_rom_13__1_), .R(_225__bF_buf4), .S(vdd) );
DFFSR DFFSR_235 ( .CLK(clk2_clkout_bF_buf17), .D(asr2_rom_12__2_), .Q(asr2_rom_13__2_), .R(_225__bF_buf3), .S(vdd) );
DFFSR DFFSR_236 ( .CLK(clk2_clkout_bF_buf16), .D(asr2_rom_12__3_), .Q(asr2_rom_13__3_), .R(_225__bF_buf2), .S(vdd) );
DFFSR DFFSR_237 ( .CLK(clk2_clkout_bF_buf15), .D(asr2_rom_12__4_), .Q(asr2_rom_13__4_), .R(_225__bF_buf1), .S(vdd) );
DFFSR DFFSR_238 ( .CLK(clk2_clkout_bF_buf14), .D(asr2_rom_12__5_), .Q(asr2_rom_13__5_), .R(_225__bF_buf0), .S(vdd) );
DFFSR DFFSR_239 ( .CLK(clk2_clkout_bF_buf13), .D(asr2_rom_12__6_), .Q(asr2_rom_13__6_), .R(_225__bF_buf10), .S(vdd) );
DFFSR DFFSR_240 ( .CLK(clk2_clkout_bF_buf12), .D(asr2_rom_12__7_), .Q(asr2_rom_13__7_), .R(_225__bF_buf9), .S(vdd) );
DFFSR DFFSR_241 ( .CLK(clk2_clkout_bF_buf11), .D(asr2_rom_13__0_), .Q(asr2_rom_14__0_), .R(_225__bF_buf8), .S(vdd) );
DFFSR DFFSR_242 ( .CLK(clk2_clkout_bF_buf10), .D(asr2_rom_13__1_), .Q(asr2_rom_14__1_), .R(_225__bF_buf7), .S(vdd) );
DFFSR DFFSR_243 ( .CLK(clk2_clkout_bF_buf9), .D(asr2_rom_13__2_), .Q(asr2_rom_14__2_), .R(_225__bF_buf6), .S(vdd) );
DFFSR DFFSR_244 ( .CLK(clk2_clkout_bF_buf8), .D(asr2_rom_13__3_), .Q(asr2_rom_14__3_), .R(_225__bF_buf5), .S(vdd) );
DFFSR DFFSR_245 ( .CLK(clk2_clkout_bF_buf7), .D(asr2_rom_13__4_), .Q(asr2_rom_14__4_), .R(_225__bF_buf4), .S(vdd) );
DFFSR DFFSR_246 ( .CLK(clk2_clkout_bF_buf6), .D(asr2_rom_13__5_), .Q(asr2_rom_14__5_), .R(_225__bF_buf3), .S(vdd) );
DFFSR DFFSR_247 ( .CLK(clk2_clkout_bF_buf5), .D(asr2_rom_13__6_), .Q(asr2_rom_14__6_), .R(_225__bF_buf2), .S(vdd) );
DFFSR DFFSR_248 ( .CLK(clk2_clkout_bF_buf4), .D(asr2_rom_13__7_), .Q(asr2_rom_14__7_), .R(_225__bF_buf1), .S(vdd) );
DFFSR DFFSR_249 ( .CLK(clk2_clkout_bF_buf3), .D(asr2_rom_14__0_), .Q(asr2_en_0_), .R(_225__bF_buf0), .S(vdd) );
DFFSR DFFSR_250 ( .CLK(clk2_clkout_bF_buf2), .D(asr2_rom_14__1_), .Q(asr2_en_1_), .R(_225__bF_buf10), .S(vdd) );
DFFSR DFFSR_251 ( .CLK(clk2_clkout_bF_buf1), .D(asr2_rom_14__2_), .Q(asr2_en_2_), .R(_225__bF_buf9), .S(vdd) );
DFFSR DFFSR_252 ( .CLK(clk2_clkout_bF_buf0), .D(asr2_rom_14__3_), .Q(asr2_en_3_), .R(_225__bF_buf8), .S(vdd) );
DFFSR DFFSR_253 ( .CLK(clk2_clkout_bF_buf41), .D(asr2_rom_14__4_), .Q(asr2_en_4_), .R(_225__bF_buf7), .S(vdd) );
DFFSR DFFSR_254 ( .CLK(clk2_clkout_bF_buf40), .D(asr2_rom_14__5_), .Q(asr2_en_5_), .R(_225__bF_buf6), .S(vdd) );
DFFSR DFFSR_255 ( .CLK(clk2_clkout_bF_buf39), .D(asr2_rom_14__6_), .Q(asr2_en_6_), .R(_225__bF_buf5), .S(vdd) );
DFFSR DFFSR_256 ( .CLK(clk2_clkout_bF_buf38), .D(asr2_rom_14__7_), .Q(asr2_en_7_), .R(_225__bF_buf4), .S(vdd) );
NOR2X1 NOR2X1_59 ( .A(rst_bF_buf3), .B(clk2_div_0_), .Y(_451__0_) );
INVX1 INVX1_119 ( .A(rst_bF_buf2), .Y(_452_) );
OAI21X1 OAI21X1_17 ( .A(clk2_div_0_), .B(clk2_div_1_), .C(_452_), .Y(_453_) );
AOI21X1 AOI21X1_1 ( .A(clk2_div_0_), .B(clk2_div_1_), .C(_453_), .Y(_451__1_) );
NAND3X1 NAND3X1_129 ( .A(clk2_div_0_), .B(clk2_div_1_), .C(clk2_div_2_), .Y(_454_) );
INVX1 INVX1_120 ( .A(clk2_div_2_), .Y(_455_) );
NAND2X1 NAND2X1_53 ( .A(clk2_div_0_), .B(clk2_div_1_), .Y(_456_) );
AOI21X1 AOI21X1_2 ( .A(_456_), .B(_455_), .C(rst_bF_buf1), .Y(_457_) );
AND2X2 AND2X2_27 ( .A(_457_), .B(_454_), .Y(_451__2_) );
AOI21X1 AOI21X1_3 ( .A(_454_), .B(clk2_clkout_bF_buf37), .C(rst_bF_buf0), .Y(_458_) );
OAI21X1 OAI21X1_18 ( .A(clk2_clkout_bF_buf36), .B(_454_), .C(_458_), .Y(_450_) );
DFFPOSX1 DFFPOSX1_1 ( .CLK(clk_bF_buf6), .D(_450_), .Q(clk2_clkout) );
DFFPOSX1 DFFPOSX1_2 ( .CLK(clk_bF_buf5), .D(_451__0_), .Q(clk2_div_0_) );
DFFPOSX1 DFFPOSX1_3 ( .CLK(clk_bF_buf4), .D(_451__1_), .Q(clk2_div_1_) );
DFFPOSX1 DFFPOSX1_4 ( .CLK(clk_bF_buf3), .D(_451__2_), .Q(clk2_div_2_) );
OR2X2 OR2X2_1 ( .A(counterup_counter_1_), .B(counterup_counter_0_bF_buf0_), .Y(_462_) );
INVX1 INVX1_121 ( .A(counterup_counter_3_), .Y(_463_) );
INVX1 INVX1_122 ( .A(counterup_counter_2_), .Y(_464_) );
INVX1 INVX1_123 ( .A(rst_bF_buf5), .Y(_460_) );
NAND3X1 NAND3X1_130 ( .A(_463_), .B(_464_), .C(_460_), .Y(_461_) );
NOR2X1 NOR2X1_60 ( .A(_462_), .B(_461_), .Y(_459_) );
DFFPOSX1 DFFPOSX1_5 ( .CLK(clk_bF_buf2), .D(_459_), .Q(comp_dataout) );
INVX1 INVX1_124 ( .A(rst_bF_buf4), .Y(_466_) );
NAND2X1 NAND2X1_54 ( .A(counterdown_counter_0_), .B(_466_), .Y(_465__0_) );
AOI21X1 AOI21X1_4 ( .A(counterdown_counter_0_), .B(counterdown_counter_1_), .C(rst_bF_buf3), .Y(_467_) );
OAI21X1 OAI21X1_19 ( .A(counterdown_counter_0_), .B(counterdown_counter_1_), .C(_467_), .Y(_465__1_) );
INVX1 INVX1_125 ( .A(counterdown_counter_0_), .Y(_468_) );
INVX1 INVX1_126 ( .A(counterdown_counter_1_), .Y(_469_) );
INVX1 INVX1_127 ( .A(counterdown_counter_2_), .Y(_470_) );
NAND3X1 NAND3X1_131 ( .A(_468_), .B(_469_), .C(_470_), .Y(_471_) );
OAI21X1 OAI21X1_20 ( .A(counterdown_counter_0_), .B(counterdown_counter_1_), .C(counterdown_counter_2_), .Y(_472_) );
NAND3X1 NAND3X1_132 ( .A(_466_), .B(_472_), .C(_471_), .Y(_465__2_) );
NAND2X1 NAND2X1_55 ( .A(counterdown_counter_3_), .B(_471_), .Y(_473_) );
INVX1 INVX1_128 ( .A(counterdown_counter_3_), .Y(_474_) );
NOR2X1 NOR2X1_61 ( .A(counterdown_counter_0_), .B(counterdown_counter_1_), .Y(_475_) );
NAND3X1 NAND3X1_133 ( .A(_470_), .B(_474_), .C(_475_), .Y(_476_) );
NAND3X1 NAND3X1_134 ( .A(_466_), .B(_476_), .C(_473_), .Y(_465__3_) );
DFFPOSX1 DFFPOSX1_6 ( .CLK(clk_bF_buf1), .D(_465__0_), .Q(counterdown_counter_0_) );
DFFPOSX1 DFFPOSX1_7 ( .CLK(clk_bF_buf0), .D(_465__1_), .Q(counterdown_counter_1_) );
DFFPOSX1 DFFPOSX1_8 ( .CLK(clk_bF_buf6), .D(_465__2_), .Q(counterdown_counter_2_) );
DFFPOSX1 DFFPOSX1_9 ( .CLK(clk_bF_buf5), .D(_465__3_), .Q(counterdown_counter_3_) );
NOR2X1 NOR2X1_62 ( .A(counterup_counter_0_bF_buf3_), .B(rst_bF_buf2), .Y(_477__0_) );
AND2X2 AND2X2_28 ( .A(counterup_counter_0_bF_buf2_), .B(counterup_counter_1_), .Y(_478_) );
INVX1 INVX1_129 ( .A(rst_bF_buf1), .Y(_479_) );
OAI21X1 OAI21X1_21 ( .A(counterup_counter_0_bF_buf1_), .B(counterup_counter_1_), .C(_479_), .Y(_480_) );
NOR2X1 NOR2X1_63 ( .A(_478_), .B(_480_), .Y(_477__1_) );
AOI21X1 AOI21X1_5 ( .A(counterup_counter_0_bF_buf0_), .B(counterup_counter_1_), .C(counterup_counter_2_), .Y(_481_) );
NAND3X1 NAND3X1_135 ( .A(counterup_counter_0_bF_buf3_), .B(counterup_counter_1_), .C(counterup_counter_2_), .Y(_482_) );
NAND2X1 NAND2X1_56 ( .A(_479_), .B(_482_), .Y(_483_) );
NOR2X1 NOR2X1_64 ( .A(_481_), .B(_483_), .Y(_477__2_) );
NAND2X1 NAND2X1_57 ( .A(counterup_counter_3_), .B(_482_), .Y(_484_) );
INVX1 INVX1_130 ( .A(counterup_counter_3_), .Y(_485_) );
NAND3X1 NAND3X1_136 ( .A(counterup_counter_2_), .B(_485_), .C(_478_), .Y(_486_) );
AOI21X1 AOI21X1_6 ( .A(_486_), .B(_484_), .C(rst_bF_buf0), .Y(_477__3_) );
DFFPOSX1 DFFPOSX1_10 ( .CLK(clk_bF_buf4), .D(_477__0_), .Q(counterup_counter_0_) );
DFFPOSX1 DFFPOSX1_11 ( .CLK(clk_bF_buf3), .D(_477__1_), .Q(counterup_counter_1_) );
DFFPOSX1 DFFPOSX1_12 ( .CLK(clk_bF_buf2), .D(_477__2_), .Q(counterup_counter_2_) );
DFFPOSX1 DFFPOSX1_13 ( .CLK(clk_bF_buf1), .D(_477__3_), .Q(counterup_counter_3_) );
NAND2X1 NAND2X1_58 ( .A(rom1_data_0_bF_buf3_), .B(sumador_res_0_), .Y(_734_) );
INVX1 INVX1_131 ( .A(mac1_reset_bF_buf3), .Y(_745_) );
NAND2X1 NAND2X1_59 ( .A(mac1_dataout_0_), .B(_745_), .Y(_756_) );
XOR2X1 XOR2X1_1 ( .A(_756_), .B(_734_), .Y(_487__0_) );
INVX1 INVX1_132 ( .A(rom1_data_0_bF_buf2_), .Y(_777_) );
INVX1 INVX1_133 ( .A(sumador_res_0_), .Y(_788_) );
INVX1 INVX1_134 ( .A(sumador_res_1_), .Y(_795_) );
INVX1 INVX1_135 ( .A(rom1_data_1_), .Y(_796_) );
OAI22X1 OAI22X1_49 ( .A(_777_), .B(_795_), .C(_788_), .D(_796_), .Y(_797_) );
NAND2X1 NAND2X1_60 ( .A(sumador_res_1_), .B(rom1_data_1_), .Y(_798_) );
OAI21X1 OAI21X1_22 ( .A(_734_), .B(_798_), .C(_797_), .Y(_799_) );
NAND3X1 NAND3X1_137 ( .A(rom1_data_0_bF_buf1_), .B(sumador_res_0_), .C(mac1_dataout_0_), .Y(_800_) );
INVX1 INVX1_136 ( .A(_800_), .Y(_801_) );
INVX1 INVX1_137 ( .A(mac1_dataout_1_), .Y(_802_) );
XOR2X1 XOR2X1_2 ( .A(_799_), .B(_802_), .Y(_803_) );
NAND2X1 NAND2X1_61 ( .A(_801_), .B(_803_), .Y(_804_) );
OR2X2 OR2X2_2 ( .A(_803_), .B(_801_), .Y(_805_) );
NAND3X1 NAND3X1_138 ( .A(_745_), .B(_804_), .C(_805_), .Y(_806_) );
OAI21X1 OAI21X1_23 ( .A(_745_), .B(_799_), .C(_806_), .Y(_487__1_) );
NAND2X1 NAND2X1_62 ( .A(sumador_res_0_), .B(rom1_data_2_), .Y(_807_) );
INVX1 INVX1_138 ( .A(_807_), .Y(_808_) );
AND2X2 AND2X2_29 ( .A(rom1_data_0_bF_buf0_), .B(sumador_res_2_), .Y(_809_) );
NAND3X1 NAND3X1_139 ( .A(sumador_res_1_), .B(rom1_data_1_), .C(_809_), .Y(_810_) );
AOI22X1 AOI22X1_17 ( .A(rom1_data_0_bF_buf3_), .B(sumador_res_2_), .C(sumador_res_1_), .D(rom1_data_1_), .Y(_811_) );
INVX1 INVX1_139 ( .A(_811_), .Y(_812_) );
NAND3X1 NAND3X1_140 ( .A(_812_), .B(_808_), .C(_810_), .Y(_813_) );
NAND2X1 NAND2X1_63 ( .A(rom1_data_0_bF_buf2_), .B(sumador_res_2_), .Y(_814_) );
NOR2X1 NOR2X1_65 ( .A(_798_), .B(_814_), .Y(_815_) );
OAI21X1 OAI21X1_24 ( .A(_811_), .B(_815_), .C(_807_), .Y(_816_) );
NAND2X1 NAND2X1_64 ( .A(_813_), .B(_816_), .Y(_817_) );
OAI21X1 OAI21X1_25 ( .A(_734_), .B(_798_), .C(_817_), .Y(_818_) );
NOR2X1 NOR2X1_66 ( .A(_734_), .B(_798_), .Y(_819_) );
NAND3X1 NAND3X1_141 ( .A(_819_), .B(_813_), .C(_816_), .Y(_820_) );
NAND2X1 NAND2X1_65 ( .A(_820_), .B(_818_), .Y(_821_) );
OAI21X1 OAI21X1_26 ( .A(_802_), .B(_799_), .C(_804_), .Y(_822_) );
INVX1 INVX1_140 ( .A(_822_), .Y(_823_) );
NAND3X1 NAND3X1_142 ( .A(mac1_dataout_2_), .B(_820_), .C(_818_), .Y(_824_) );
INVX1 INVX1_141 ( .A(_824_), .Y(_825_) );
AOI21X1 AOI21X1_7 ( .A(_818_), .B(_820_), .C(mac1_dataout_2_), .Y(_826_) );
NOR2X1 NOR2X1_67 ( .A(_826_), .B(_825_), .Y(_827_) );
AND2X2 AND2X2_30 ( .A(_827_), .B(_823_), .Y(_828_) );
NOR2X1 NOR2X1_68 ( .A(_823_), .B(_827_), .Y(_829_) );
OAI21X1 OAI21X1_27 ( .A(_829_), .B(_828_), .C(_745_), .Y(_830_) );
OAI21X1 OAI21X1_28 ( .A(_745_), .B(_821_), .C(_830_), .Y(_487__2_) );
OAI21X1 OAI21X1_29 ( .A(_826_), .B(_823_), .C(_824_), .Y(_831_) );
INVX1 INVX1_142 ( .A(_820_), .Y(_832_) );
NAND2X1 NAND2X1_66 ( .A(sumador_res_0_), .B(rom1_data_3_), .Y(_833_) );
INVX1 INVX1_143 ( .A(_833_), .Y(_834_) );
OAI21X1 OAI21X1_30 ( .A(_807_), .B(_811_), .C(_810_), .Y(_835_) );
NAND2X1 NAND2X1_67 ( .A(sumador_res_1_), .B(rom1_data_2_), .Y(_836_) );
INVX1 INVX1_144 ( .A(_836_), .Y(_837_) );
AND2X2 AND2X2_31 ( .A(rom1_data_1_), .B(sumador_res_2_), .Y(_838_) );
AND2X2 AND2X2_32 ( .A(rom1_data_0_bF_buf1_), .B(sumador_res_3_), .Y(_839_) );
NAND2X1 NAND2X1_68 ( .A(_838_), .B(_839_), .Y(_840_) );
INVX1 INVX1_145 ( .A(sumador_res_2_), .Y(_841_) );
NAND2X1 NAND2X1_69 ( .A(rom1_data_0_bF_buf0_), .B(sumador_res_3_), .Y(_842_) );
OAI21X1 OAI21X1_31 ( .A(_796_), .B(_841_), .C(_842_), .Y(_843_) );
NAND3X1 NAND3X1_143 ( .A(_843_), .B(_837_), .C(_840_), .Y(_844_) );
OAI21X1 OAI21X1_32 ( .A(_796_), .B(_841_), .C(_839_), .Y(_845_) );
INVX1 INVX1_146 ( .A(sumador_res_3_), .Y(_846_) );
OAI21X1 OAI21X1_33 ( .A(_777_), .B(_846_), .C(_838_), .Y(_847_) );
NAND3X1 NAND3X1_144 ( .A(_836_), .B(_845_), .C(_847_), .Y(_848_) );
NAND3X1 NAND3X1_145 ( .A(_844_), .B(_835_), .C(_848_), .Y(_849_) );
AOI21X1 AOI21X1_8 ( .A(_808_), .B(_812_), .C(_815_), .Y(_850_) );
NAND3X1 NAND3X1_146 ( .A(_836_), .B(_843_), .C(_840_), .Y(_851_) );
NAND3X1 NAND3X1_147 ( .A(_837_), .B(_845_), .C(_847_), .Y(_852_) );
NAND3X1 NAND3X1_148 ( .A(_851_), .B(_852_), .C(_850_), .Y(_488_) );
NAND3X1 NAND3X1_149 ( .A(_834_), .B(_849_), .C(_488_), .Y(_489_) );
NAND3X1 NAND3X1_150 ( .A(_844_), .B(_848_), .C(_850_), .Y(_490_) );
NAND3X1 NAND3X1_151 ( .A(_851_), .B(_835_), .C(_852_), .Y(_491_) );
NAND3X1 NAND3X1_152 ( .A(_833_), .B(_491_), .C(_490_), .Y(_492_) );
AOI21X1 AOI21X1_9 ( .A(_489_), .B(_492_), .C(_832_), .Y(_493_) );
INVX1 INVX1_147 ( .A(_493_), .Y(_494_) );
NAND3X1 NAND3X1_153 ( .A(_832_), .B(_489_), .C(_492_), .Y(_495_) );
NAND3X1 NAND3X1_154 ( .A(mac1_dataout_3_), .B(_495_), .C(_494_), .Y(_496_) );
INVX1 INVX1_148 ( .A(mac1_dataout_3_), .Y(_497_) );
INVX1 INVX1_149 ( .A(_495_), .Y(_498_) );
OAI21X1 OAI21X1_34 ( .A(_493_), .B(_498_), .C(_497_), .Y(_499_) );
NAND2X1 NAND2X1_70 ( .A(_496_), .B(_499_), .Y(_500_) );
XOR2X1 XOR2X1_3 ( .A(_500_), .B(_831_), .Y(_501_) );
NAND3X1 NAND3X1_155 ( .A(mac1_reset_bF_buf2), .B(_495_), .C(_494_), .Y(_502_) );
OAI21X1 OAI21X1_35 ( .A(mac1_reset_bF_buf1), .B(_501_), .C(_502_), .Y(_487__3_) );
NAND2X1 NAND2X1_71 ( .A(sumador_res_1_), .B(rom1_data_4_), .Y(_503_) );
INVX1 INVX1_150 ( .A(rom1_data_4_), .Y(_504_) );
NAND2X1 NAND2X1_72 ( .A(sumador_res_1_), .B(rom1_data_3_), .Y(_505_) );
OAI21X1 OAI21X1_36 ( .A(_788_), .B(_504_), .C(_505_), .Y(_506_) );
OAI21X1 OAI21X1_37 ( .A(_833_), .B(_503_), .C(_506_), .Y(_507_) );
AOI22X1 AOI22X1_18 ( .A(rom1_data_0_bF_buf3_), .B(sumador_res_3_), .C(rom1_data_1_), .D(sumador_res_2_), .Y(_508_) );
OAI21X1 OAI21X1_38 ( .A(_836_), .B(_508_), .C(_840_), .Y(_509_) );
NAND2X1 NAND2X1_73 ( .A(sumador_res_2_), .B(rom1_data_2_), .Y(_510_) );
INVX1 INVX1_151 ( .A(_510_), .Y(_511_) );
AND2X2 AND2X2_33 ( .A(rom1_data_1_), .B(sumador_res_4_), .Y(_512_) );
NAND2X1 NAND2X1_74 ( .A(_839_), .B(_512_), .Y(_513_) );
NAND2X1 NAND2X1_75 ( .A(rom1_data_1_), .B(sumador_res_3_), .Y(_514_) );
NAND2X1 NAND2X1_76 ( .A(rom1_data_0_bF_buf2_), .B(sumador_res_4_), .Y(_515_) );
NAND2X1 NAND2X1_77 ( .A(_514_), .B(_515_), .Y(_516_) );
NAND3X1 NAND3X1_156 ( .A(_511_), .B(_516_), .C(_513_), .Y(_517_) );
NAND3X1 NAND3X1_157 ( .A(rom1_data_0_bF_buf1_), .B(sumador_res_4_), .C(_514_), .Y(_518_) );
AND2X2 AND2X2_34 ( .A(rom1_data_1_), .B(sumador_res_3_), .Y(_519_) );
NAND2X1 NAND2X1_78 ( .A(_515_), .B(_519_), .Y(_520_) );
NAND3X1 NAND3X1_158 ( .A(_510_), .B(_518_), .C(_520_), .Y(_521_) );
NAND3X1 NAND3X1_159 ( .A(_509_), .B(_517_), .C(_521_), .Y(_522_) );
AOI22X1 AOI22X1_19 ( .A(_809_), .B(_519_), .C(_843_), .D(_837_), .Y(_523_) );
NAND3X1 NAND3X1_160 ( .A(_510_), .B(_516_), .C(_513_), .Y(_524_) );
NAND3X1 NAND3X1_161 ( .A(_511_), .B(_518_), .C(_520_), .Y(_525_) );
NAND3X1 NAND3X1_162 ( .A(_525_), .B(_524_), .C(_523_), .Y(_526_) );
NAND3X1 NAND3X1_163 ( .A(_507_), .B(_522_), .C(_526_), .Y(_527_) );
INVX1 INVX1_152 ( .A(_507_), .Y(_528_) );
AOI21X1 AOI21X1_10 ( .A(_524_), .B(_525_), .C(_523_), .Y(_529_) );
AOI21X1 AOI21X1_11 ( .A(_517_), .B(_521_), .C(_509_), .Y(_530_) );
OAI21X1 OAI21X1_39 ( .A(_530_), .B(_529_), .C(_528_), .Y(_531_) );
AOI22X1 AOI22X1_20 ( .A(_849_), .B(_489_), .C(_531_), .D(_527_), .Y(_532_) );
AOI21X1 AOI21X1_12 ( .A(_848_), .B(_844_), .C(_835_), .Y(_533_) );
OAI21X1 OAI21X1_40 ( .A(_833_), .B(_533_), .C(_849_), .Y(_534_) );
NAND3X1 NAND3X1_164 ( .A(_528_), .B(_522_), .C(_526_), .Y(_535_) );
OAI21X1 OAI21X1_41 ( .A(_530_), .B(_529_), .C(_507_), .Y(_536_) );
AOI21X1 AOI21X1_13 ( .A(_535_), .B(_536_), .C(_534_), .Y(_537_) );
OAI21X1 OAI21X1_42 ( .A(_532_), .B(_537_), .C(_495_), .Y(_538_) );
NAND3X1 NAND3X1_165 ( .A(_535_), .B(_536_), .C(_534_), .Y(_539_) );
AOI21X1 AOI21X1_14 ( .A(_851_), .B(_852_), .C(_850_), .Y(_540_) );
AOI21X1 AOI21X1_15 ( .A(_834_), .B(_488_), .C(_540_), .Y(_541_) );
NAND3X1 NAND3X1_166 ( .A(_527_), .B(_531_), .C(_541_), .Y(_542_) );
NAND3X1 NAND3X1_167 ( .A(_539_), .B(_542_), .C(_498_), .Y(_543_) );
NAND2X1 NAND2X1_79 ( .A(_538_), .B(_543_), .Y(_544_) );
INVX1 INVX1_153 ( .A(_826_), .Y(_545_) );
AOI21X1 AOI21X1_16 ( .A(_545_), .B(_822_), .C(_825_), .Y(_546_) );
AOI21X1 AOI21X1_17 ( .A(_494_), .B(_495_), .C(mac1_dataout_3_), .Y(_547_) );
OAI21X1 OAI21X1_43 ( .A(_546_), .B(_547_), .C(_496_), .Y(_548_) );
NAND3X1 NAND3X1_168 ( .A(mac1_dataout_4_), .B(_538_), .C(_543_), .Y(_549_) );
INVX1 INVX1_154 ( .A(mac1_dataout_4_), .Y(_550_) );
NAND2X1 NAND2X1_80 ( .A(_550_), .B(_544_), .Y(_551_) );
NAND3X1 NAND3X1_169 ( .A(_549_), .B(_548_), .C(_551_), .Y(_552_) );
INVX1 INVX1_155 ( .A(_496_), .Y(_553_) );
AOI21X1 AOI21X1_18 ( .A(_499_), .B(_831_), .C(_553_), .Y(_554_) );
INVX1 INVX1_156 ( .A(_549_), .Y(_555_) );
AOI21X1 AOI21X1_19 ( .A(_543_), .B(_538_), .C(mac1_dataout_4_), .Y(_556_) );
OAI21X1 OAI21X1_44 ( .A(_556_), .B(_555_), .C(_554_), .Y(_557_) );
NAND3X1 NAND3X1_170 ( .A(_745_), .B(_552_), .C(_557_), .Y(_558_) );
OAI21X1 OAI21X1_45 ( .A(_745_), .B(_544_), .C(_558_), .Y(_487__4_) );
NOR3X1 NOR3X1_5 ( .A(_495_), .B(_532_), .C(_537_), .Y(_559_) );
AND2X2 AND2X2_35 ( .A(sumador_res_1_), .B(rom1_data_4_), .Y(_560_) );
NAND2X1 NAND2X1_81 ( .A(_560_), .B(_834_), .Y(_561_) );
INVX1 INVX1_157 ( .A(_561_), .Y(_562_) );
OAI21X1 OAI21X1_46 ( .A(_507_), .B(_530_), .C(_522_), .Y(_563_) );
NAND2X1 NAND2X1_82 ( .A(sumador_res_0_), .B(gnd), .Y(_564_) );
INVX1 INVX1_158 ( .A(_564_), .Y(_565_) );
AND2X2 AND2X2_36 ( .A(sumador_res_2_), .B(rom1_data_3_), .Y(_566_) );
NAND2X1 NAND2X1_83 ( .A(_560_), .B(_566_), .Y(_567_) );
INVX1 INVX1_159 ( .A(rom1_data_3_), .Y(_568_) );
OAI21X1 OAI21X1_47 ( .A(_841_), .B(_568_), .C(_503_), .Y(_569_) );
NAND3X1 NAND3X1_171 ( .A(_569_), .B(_565_), .C(_567_), .Y(_570_) );
OAI21X1 OAI21X1_48 ( .A(_795_), .B(_504_), .C(_566_), .Y(_571_) );
OAI21X1 OAI21X1_49 ( .A(_841_), .B(_568_), .C(_560_), .Y(_572_) );
NAND3X1 NAND3X1_172 ( .A(_564_), .B(_571_), .C(_572_), .Y(_573_) );
AOI22X1 AOI22X1_21 ( .A(_839_), .B(_512_), .C(_516_), .D(_511_), .Y(_574_) );
NAND2X1 NAND2X1_84 ( .A(rom1_data_2_), .B(sumador_res_3_), .Y(_575_) );
INVX1 INVX1_160 ( .A(_575_), .Y(_576_) );
AND2X2 AND2X2_37 ( .A(rom1_data_0_bF_buf0_), .B(sumador_res_5_), .Y(_577_) );
NAND2X1 NAND2X1_85 ( .A(_512_), .B(_577_), .Y(_578_) );
INVX1 INVX1_161 ( .A(sumador_res_5_), .Y(_579_) );
NAND2X1 NAND2X1_86 ( .A(rom1_data_1_), .B(sumador_res_4_), .Y(_580_) );
OAI21X1 OAI21X1_50 ( .A(_777_), .B(_579_), .C(_580_), .Y(_581_) );
NAND3X1 NAND3X1_173 ( .A(_576_), .B(_581_), .C(_578_), .Y(_582_) );
NAND3X1 NAND3X1_174 ( .A(rom1_data_0_bF_buf3_), .B(sumador_res_5_), .C(_580_), .Y(_583_) );
NAND2X1 NAND2X1_87 ( .A(rom1_data_0_bF_buf2_), .B(sumador_res_5_), .Y(_584_) );
NAND3X1 NAND3X1_175 ( .A(rom1_data_1_), .B(sumador_res_4_), .C(_584_), .Y(_585_) );
NAND3X1 NAND3X1_176 ( .A(_575_), .B(_583_), .C(_585_), .Y(_586_) );
NAND3X1 NAND3X1_177 ( .A(_574_), .B(_586_), .C(_582_), .Y(_587_) );
AOI22X1 AOI22X1_22 ( .A(rom1_data_0_bF_buf1_), .B(sumador_res_4_), .C(rom1_data_1_), .D(sumador_res_3_), .Y(_588_) );
OAI22X1 OAI22X1_50 ( .A(_842_), .B(_580_), .C(_510_), .D(_588_), .Y(_589_) );
NAND3X1 NAND3X1_178 ( .A(_575_), .B(_581_), .C(_578_), .Y(_590_) );
NAND3X1 NAND3X1_179 ( .A(_576_), .B(_583_), .C(_585_), .Y(_591_) );
NAND3X1 NAND3X1_180 ( .A(_589_), .B(_591_), .C(_590_), .Y(_592_) );
AOI22X1 AOI22X1_23 ( .A(_570_), .B(_573_), .C(_587_), .D(_592_), .Y(_593_) );
NAND3X1 NAND3X1_181 ( .A(_564_), .B(_569_), .C(_567_), .Y(_594_) );
NAND3X1 NAND3X1_182 ( .A(_565_), .B(_571_), .C(_572_), .Y(_595_) );
NAND3X1 NAND3X1_183 ( .A(_589_), .B(_586_), .C(_582_), .Y(_596_) );
NAND3X1 NAND3X1_184 ( .A(_574_), .B(_591_), .C(_590_), .Y(_597_) );
AOI22X1 AOI22X1_24 ( .A(_594_), .B(_595_), .C(_596_), .D(_597_), .Y(_598_) );
OAI21X1 OAI21X1_51 ( .A(_593_), .B(_598_), .C(_563_), .Y(_599_) );
AOI21X1 AOI21X1_20 ( .A(_528_), .B(_526_), .C(_529_), .Y(_600_) );
NAND2X1 NAND2X1_88 ( .A(_570_), .B(_573_), .Y(_601_) );
AOI21X1 AOI21X1_21 ( .A(_587_), .B(_592_), .C(_601_), .Y(_602_) );
NAND2X1 NAND2X1_89 ( .A(_594_), .B(_595_), .Y(_603_) );
AOI21X1 AOI21X1_22 ( .A(_596_), .B(_597_), .C(_603_), .Y(_604_) );
OAI21X1 OAI21X1_52 ( .A(_604_), .B(_602_), .C(_600_), .Y(_605_) );
NAND3X1 NAND3X1_185 ( .A(_562_), .B(_599_), .C(_605_), .Y(_606_) );
OAI21X1 OAI21X1_53 ( .A(_593_), .B(_598_), .C(_600_), .Y(_607_) );
OAI21X1 OAI21X1_54 ( .A(_604_), .B(_602_), .C(_563_), .Y(_608_) );
NAND3X1 NAND3X1_186 ( .A(_561_), .B(_607_), .C(_608_), .Y(_609_) );
NAND3X1 NAND3X1_187 ( .A(_532_), .B(_606_), .C(_609_), .Y(_610_) );
NAND3X1 NAND3X1_188 ( .A(_561_), .B(_599_), .C(_605_), .Y(_611_) );
NAND3X1 NAND3X1_189 ( .A(_562_), .B(_607_), .C(_608_), .Y(_612_) );
NAND3X1 NAND3X1_190 ( .A(_539_), .B(_611_), .C(_612_), .Y(_613_) );
NAND3X1 NAND3X1_191 ( .A(_559_), .B(_610_), .C(_613_), .Y(_614_) );
NAND3X1 NAND3X1_192 ( .A(_539_), .B(_606_), .C(_609_), .Y(_615_) );
NAND3X1 NAND3X1_193 ( .A(_532_), .B(_611_), .C(_612_), .Y(_616_) );
NAND3X1 NAND3X1_194 ( .A(_543_), .B(_615_), .C(_616_), .Y(_617_) );
NAND2X1 NAND2X1_90 ( .A(_614_), .B(_617_), .Y(_618_) );
OAI21X1 OAI21X1_55 ( .A(_556_), .B(_554_), .C(_549_), .Y(_619_) );
NAND3X1 NAND3X1_195 ( .A(mac1_dataout_5_), .B(_614_), .C(_617_), .Y(_620_) );
INVX1 INVX1_162 ( .A(mac1_dataout_5_), .Y(_621_) );
NAND2X1 NAND2X1_91 ( .A(_621_), .B(_618_), .Y(_622_) );
NAND3X1 NAND3X1_196 ( .A(_620_), .B(_622_), .C(_619_), .Y(_623_) );
AOI21X1 AOI21X1_23 ( .A(_548_), .B(_551_), .C(_555_), .Y(_624_) );
INVX1 INVX1_163 ( .A(_620_), .Y(_625_) );
AOI21X1 AOI21X1_24 ( .A(_614_), .B(_617_), .C(mac1_dataout_5_), .Y(_626_) );
OAI21X1 OAI21X1_56 ( .A(_626_), .B(_625_), .C(_624_), .Y(_627_) );
NAND3X1 NAND3X1_197 ( .A(_745_), .B(_623_), .C(_627_), .Y(_628_) );
OAI21X1 OAI21X1_57 ( .A(_745_), .B(_618_), .C(_628_), .Y(_487__5_) );
AOI21X1 AOI21X1_25 ( .A(_615_), .B(_616_), .C(_543_), .Y(_629_) );
AOI21X1 AOI21X1_26 ( .A(_612_), .B(_611_), .C(_539_), .Y(_630_) );
NAND3X1 NAND3X1_198 ( .A(_596_), .B(_597_), .C(_603_), .Y(_631_) );
AOI21X1 AOI21X1_27 ( .A(_590_), .B(_591_), .C(_574_), .Y(_632_) );
AOI21X1 AOI21X1_28 ( .A(_582_), .B(_586_), .C(_589_), .Y(_633_) );
OAI21X1 OAI21X1_58 ( .A(_632_), .B(_633_), .C(_601_), .Y(_634_) );
AOI21X1 AOI21X1_29 ( .A(_634_), .B(_631_), .C(_563_), .Y(_635_) );
OAI21X1 OAI21X1_59 ( .A(_561_), .B(_635_), .C(_599_), .Y(_636_) );
AND2X2 AND2X2_38 ( .A(sumador_res_0_), .B(gnd), .Y(_637_) );
NAND2X1 NAND2X1_92 ( .A(sumador_res_2_), .B(rom1_data_4_), .Y(_638_) );
OAI21X1 OAI21X1_60 ( .A(_505_), .B(_638_), .C(_570_), .Y(_639_) );
XNOR2X1 XNOR2X1_1 ( .A(_639_), .B(_637_), .Y(_640_) );
INVX1 INVX1_164 ( .A(_640_), .Y(_641_) );
OAI21X1 OAI21X1_61 ( .A(_601_), .B(_633_), .C(_596_), .Y(_642_) );
INVX1 INVX1_165 ( .A(gnd), .Y(_643_) );
NOR2X1 NOR2X1_69 ( .A(_795_), .B(_643_), .Y(_644_) );
NAND2X1 NAND2X1_93 ( .A(sumador_res_3_), .B(rom1_data_3_), .Y(_645_) );
XOR2X1 XOR2X1_4 ( .A(_638_), .B(_645_), .Y(_646_) );
NAND2X1 NAND2X1_94 ( .A(_644_), .B(_646_), .Y(_647_) );
INVX1 INVX1_166 ( .A(_566_), .Y(_648_) );
NAND2X1 NAND2X1_95 ( .A(sumador_res_3_), .B(rom1_data_4_), .Y(_649_) );
OAI21X1 OAI21X1_62 ( .A(_846_), .B(_568_), .C(_638_), .Y(_650_) );
OAI21X1 OAI21X1_63 ( .A(_649_), .B(_648_), .C(_650_), .Y(_651_) );
OAI21X1 OAI21X1_64 ( .A(_795_), .B(_643_), .C(_651_), .Y(_652_) );
NOR2X1 NOR2X1_70 ( .A(_580_), .B(_584_), .Y(_653_) );
AOI21X1 AOI21X1_30 ( .A(_576_), .B(_581_), .C(_653_), .Y(_654_) );
NAND2X1 NAND2X1_96 ( .A(rom1_data_2_), .B(sumador_res_4_), .Y(_655_) );
INVX1 INVX1_167 ( .A(_655_), .Y(_656_) );
NAND3X1 NAND3X1_199 ( .A(rom1_data_1_), .B(sumador_res_6_), .C(_577_), .Y(_657_) );
AOI22X1 AOI22X1_25 ( .A(rom1_data_0_bF_buf0_), .B(sumador_res_6_), .C(rom1_data_1_), .D(sumador_res_5_), .Y(_658_) );
INVX1 INVX1_168 ( .A(_658_), .Y(_659_) );
NAND3X1 NAND3X1_200 ( .A(_659_), .B(_656_), .C(_657_), .Y(_660_) );
NAND2X1 NAND2X1_97 ( .A(rom1_data_1_), .B(sumador_res_6_), .Y(_661_) );
NOR2X1 NOR2X1_71 ( .A(_584_), .B(_661_), .Y(_662_) );
OAI21X1 OAI21X1_65 ( .A(_658_), .B(_662_), .C(_655_), .Y(_663_) );
NAND3X1 NAND3X1_201 ( .A(_660_), .B(_663_), .C(_654_), .Y(_664_) );
AND2X2 AND2X2_39 ( .A(_580_), .B(_584_), .Y(_665_) );
OAI21X1 OAI21X1_66 ( .A(_575_), .B(_665_), .C(_578_), .Y(_666_) );
NAND3X1 NAND3X1_202 ( .A(_655_), .B(_659_), .C(_657_), .Y(_667_) );
OAI21X1 OAI21X1_67 ( .A(_658_), .B(_662_), .C(_656_), .Y(_668_) );
NAND3X1 NAND3X1_203 ( .A(_667_), .B(_668_), .C(_666_), .Y(_669_) );
AOI22X1 AOI22X1_26 ( .A(_647_), .B(_652_), .C(_664_), .D(_669_), .Y(_670_) );
OAI21X1 OAI21X1_68 ( .A(_795_), .B(_643_), .C(_646_), .Y(_671_) );
NAND2X1 NAND2X1_98 ( .A(_644_), .B(_651_), .Y(_672_) );
NAND3X1 NAND3X1_204 ( .A(_660_), .B(_663_), .C(_666_), .Y(_673_) );
NAND3X1 NAND3X1_205 ( .A(_667_), .B(_668_), .C(_654_), .Y(_674_) );
AOI22X1 AOI22X1_27 ( .A(_671_), .B(_672_), .C(_674_), .D(_673_), .Y(_675_) );
OAI21X1 OAI21X1_69 ( .A(_670_), .B(_675_), .C(_642_), .Y(_676_) );
AOI21X1 AOI21X1_31 ( .A(_603_), .B(_597_), .C(_632_), .Y(_677_) );
AOI22X1 AOI22X1_28 ( .A(_671_), .B(_672_), .C(_664_), .D(_669_), .Y(_678_) );
AOI22X1 AOI22X1_29 ( .A(_647_), .B(_652_), .C(_674_), .D(_673_), .Y(_679_) );
OAI21X1 OAI21X1_70 ( .A(_678_), .B(_679_), .C(_677_), .Y(_680_) );
NAND3X1 NAND3X1_206 ( .A(_676_), .B(_641_), .C(_680_), .Y(_681_) );
OAI21X1 OAI21X1_71 ( .A(_670_), .B(_675_), .C(_677_), .Y(_682_) );
OAI21X1 OAI21X1_72 ( .A(_678_), .B(_679_), .C(_642_), .Y(_683_) );
NAND3X1 NAND3X1_207 ( .A(_640_), .B(_682_), .C(_683_), .Y(_684_) );
NAND3X1 NAND3X1_208 ( .A(_684_), .B(_681_), .C(_636_), .Y(_685_) );
NAND3X1 NAND3X1_209 ( .A(_596_), .B(_601_), .C(_597_), .Y(_686_) );
OAI21X1 OAI21X1_73 ( .A(_632_), .B(_633_), .C(_603_), .Y(_687_) );
AOI21X1 AOI21X1_32 ( .A(_687_), .B(_686_), .C(_600_), .Y(_688_) );
AOI21X1 AOI21X1_33 ( .A(_562_), .B(_605_), .C(_688_), .Y(_689_) );
NAND3X1 NAND3X1_210 ( .A(_640_), .B(_676_), .C(_680_), .Y(_690_) );
NAND3X1 NAND3X1_211 ( .A(_682_), .B(_641_), .C(_683_), .Y(_691_) );
NAND3X1 NAND3X1_212 ( .A(_690_), .B(_691_), .C(_689_), .Y(_692_) );
NAND3X1 NAND3X1_213 ( .A(_630_), .B(_692_), .C(_685_), .Y(_693_) );
NAND3X1 NAND3X1_214 ( .A(_684_), .B(_681_), .C(_689_), .Y(_694_) );
NAND3X1 NAND3X1_215 ( .A(_690_), .B(_691_), .C(_636_), .Y(_695_) );
NAND3X1 NAND3X1_216 ( .A(_610_), .B(_694_), .C(_695_), .Y(_696_) );
NAND3X1 NAND3X1_217 ( .A(_629_), .B(_693_), .C(_696_), .Y(_697_) );
NAND3X1 NAND3X1_218 ( .A(_610_), .B(_692_), .C(_685_), .Y(_698_) );
NAND3X1 NAND3X1_219 ( .A(_630_), .B(_694_), .C(_695_), .Y(_699_) );
NAND3X1 NAND3X1_220 ( .A(_614_), .B(_698_), .C(_699_), .Y(_700_) );
NAND2X1 NAND2X1_99 ( .A(_697_), .B(_700_), .Y(_701_) );
OAI21X1 OAI21X1_74 ( .A(_626_), .B(_624_), .C(_620_), .Y(_702_) );
NAND3X1 NAND3X1_221 ( .A(mac1_dataout_6_), .B(_697_), .C(_700_), .Y(_703_) );
INVX1 INVX1_169 ( .A(mac1_dataout_6_), .Y(_704_) );
NAND3X1 NAND3X1_222 ( .A(_614_), .B(_693_), .C(_696_), .Y(_705_) );
NAND3X1 NAND3X1_223 ( .A(_629_), .B(_698_), .C(_699_), .Y(_706_) );
NAND3X1 NAND3X1_224 ( .A(_704_), .B(_705_), .C(_706_), .Y(_707_) );
AOI21X1 AOI21X1_34 ( .A(_703_), .B(_707_), .C(_702_), .Y(_708_) );
AOI21X1 AOI21X1_35 ( .A(_619_), .B(_622_), .C(_625_), .Y(_709_) );
NAND2X1 NAND2X1_100 ( .A(_703_), .B(_707_), .Y(_710_) );
OAI21X1 OAI21X1_75 ( .A(_709_), .B(_710_), .C(_745_), .Y(_711_) );
OAI22X1 OAI22X1_51 ( .A(_745_), .B(_701_), .C(_708_), .D(_711_), .Y(_487__6_) );
NAND2X1 NAND2X1_101 ( .A(_693_), .B(_697_), .Y(_712_) );
INVX1 INVX1_170 ( .A(_712_), .Y(_713_) );
INVX1 INVX1_171 ( .A(_685_), .Y(_714_) );
NAND2X1 NAND2X1_102 ( .A(_637_), .B(_639_), .Y(_715_) );
INVX1 INVX1_172 ( .A(_715_), .Y(_716_) );
NAND2X1 NAND2X1_103 ( .A(_676_), .B(_681_), .Y(_717_) );
OAI21X1 OAI21X1_76 ( .A(_648_), .B(_649_), .C(_647_), .Y(_718_) );
NAND2X1 NAND2X1_104 ( .A(sumador_res_0_), .B(gnd), .Y(_719_) );
NAND2X1 NAND2X1_105 ( .A(sumador_res_1_), .B(gnd), .Y(_720_) );
XOR2X1 XOR2X1_5 ( .A(_719_), .B(_720_), .Y(_721_) );
XOR2X1 XOR2X1_6 ( .A(_718_), .B(_721_), .Y(_722_) );
INVX1 INVX1_173 ( .A(_722_), .Y(_723_) );
INVX1 INVX1_174 ( .A(_673_), .Y(_724_) );
OR2X2 OR2X2_3 ( .A(_678_), .B(_724_), .Y(_725_) );
INVX1 INVX1_175 ( .A(rom1_data_2_), .Y(_726_) );
NOR2X1 NOR2X1_72 ( .A(_726_), .B(_579_), .Y(_727_) );
NAND2X1 NAND2X1_106 ( .A(rom1_data_0_bF_buf3_), .B(sumador_res_7_), .Y(_728_) );
XNOR2X1 XNOR2X1_2 ( .A(_661_), .B(_728_), .Y(_729_) );
INVX1 INVX1_176 ( .A(_729_), .Y(_730_) );
NAND2X1 NAND2X1_107 ( .A(_727_), .B(_730_), .Y(_731_) );
OAI21X1 OAI21X1_77 ( .A(_726_), .B(_579_), .C(_729_), .Y(_732_) );
OAI21X1 OAI21X1_78 ( .A(_655_), .B(_658_), .C(_657_), .Y(_733_) );
INVX1 INVX1_177 ( .A(_733_), .Y(_735_) );
NAND3X1 NAND3X1_225 ( .A(_732_), .B(_735_), .C(_731_), .Y(_736_) );
NAND2X1 NAND2X1_108 ( .A(_727_), .B(_729_), .Y(_737_) );
OAI21X1 OAI21X1_79 ( .A(_726_), .B(_579_), .C(_730_), .Y(_738_) );
NAND3X1 NAND3X1_226 ( .A(_733_), .B(_737_), .C(_738_), .Y(_739_) );
NAND2X1 NAND2X1_109 ( .A(rom1_data_3_), .B(sumador_res_4_), .Y(_740_) );
XNOR2X1 XNOR2X1_3 ( .A(_649_), .B(_740_), .Y(_741_) );
NAND2X1 NAND2X1_110 ( .A(sumador_res_2_), .B(gnd), .Y(_742_) );
XOR2X1 XOR2X1_7 ( .A(_741_), .B(_742_), .Y(_743_) );
INVX1 INVX1_178 ( .A(_743_), .Y(_744_) );
NAND3X1 NAND3X1_227 ( .A(_736_), .B(_739_), .C(_744_), .Y(_746_) );
NAND3X1 NAND3X1_228 ( .A(_732_), .B(_733_), .C(_731_), .Y(_747_) );
NAND3X1 NAND3X1_229 ( .A(_735_), .B(_737_), .C(_738_), .Y(_748_) );
NAND3X1 NAND3X1_230 ( .A(_743_), .B(_747_), .C(_748_), .Y(_749_) );
NAND3X1 NAND3X1_231 ( .A(_749_), .B(_746_), .C(_725_), .Y(_750_) );
NOR2X1 NOR2X1_73 ( .A(_724_), .B(_678_), .Y(_751_) );
NAND3X1 NAND3X1_232 ( .A(_747_), .B(_748_), .C(_744_), .Y(_752_) );
NAND3X1 NAND3X1_233 ( .A(_743_), .B(_736_), .C(_739_), .Y(_753_) );
NAND3X1 NAND3X1_234 ( .A(_751_), .B(_753_), .C(_752_), .Y(_754_) );
AOI21X1 AOI21X1_36 ( .A(_750_), .B(_754_), .C(_723_), .Y(_755_) );
NAND3X1 NAND3X1_235 ( .A(_751_), .B(_749_), .C(_746_), .Y(_757_) );
NAND3X1 NAND3X1_236 ( .A(_753_), .B(_752_), .C(_725_), .Y(_758_) );
AOI21X1 AOI21X1_37 ( .A(_758_), .B(_757_), .C(_722_), .Y(_759_) );
OAI21X1 OAI21X1_80 ( .A(_755_), .B(_759_), .C(_717_), .Y(_760_) );
INVX1 INVX1_179 ( .A(_717_), .Y(_761_) );
NAND3X1 NAND3X1_237 ( .A(_722_), .B(_757_), .C(_758_), .Y(_762_) );
NAND3X1 NAND3X1_238 ( .A(_723_), .B(_754_), .C(_750_), .Y(_763_) );
NAND3X1 NAND3X1_239 ( .A(_762_), .B(_763_), .C(_761_), .Y(_764_) );
AOI21X1 AOI21X1_38 ( .A(_764_), .B(_760_), .C(_716_), .Y(_765_) );
NAND3X1 NAND3X1_240 ( .A(_717_), .B(_762_), .C(_763_), .Y(_766_) );
OAI21X1 OAI21X1_81 ( .A(_755_), .B(_759_), .C(_761_), .Y(_767_) );
AOI21X1 AOI21X1_39 ( .A(_767_), .B(_766_), .C(_715_), .Y(_768_) );
OAI21X1 OAI21X1_82 ( .A(_768_), .B(_765_), .C(_714_), .Y(_769_) );
NAND3X1 NAND3X1_241 ( .A(_715_), .B(_766_), .C(_767_), .Y(_770_) );
NAND3X1 NAND3X1_242 ( .A(_716_), .B(_760_), .C(_764_), .Y(_771_) );
NAND3X1 NAND3X1_243 ( .A(_685_), .B(_770_), .C(_771_), .Y(_772_) );
NAND3X1 NAND3X1_244 ( .A(_713_), .B(_772_), .C(_769_), .Y(_773_) );
NAND2X1 NAND2X1_111 ( .A(_760_), .B(_764_), .Y(_774_) );
XOR2X1 XOR2X1_8 ( .A(_685_), .B(_716_), .Y(_775_) );
OR2X2 OR2X2_4 ( .A(_774_), .B(_775_), .Y(_776_) );
NAND2X1 NAND2X1_112 ( .A(_775_), .B(_774_), .Y(_778_) );
NAND3X1 NAND3X1_245 ( .A(_712_), .B(_778_), .C(_776_), .Y(_779_) );
NAND2X1 NAND2X1_113 ( .A(_779_), .B(_773_), .Y(_780_) );
INVX1 INVX1_180 ( .A(mac1_dataout_7_), .Y(_781_) );
AOI21X1 AOI21X1_40 ( .A(_705_), .B(_706_), .C(_704_), .Y(_782_) );
AOI21X1 AOI21X1_41 ( .A(_702_), .B(_707_), .C(_782_), .Y(_783_) );
NAND2X1 NAND2X1_114 ( .A(_781_), .B(_783_), .Y(_784_) );
AOI21X1 AOI21X1_42 ( .A(_697_), .B(_700_), .C(mac1_dataout_6_), .Y(_785_) );
OAI21X1 OAI21X1_83 ( .A(_785_), .B(_709_), .C(_703_), .Y(_786_) );
AOI21X1 AOI21X1_43 ( .A(_786_), .B(mac1_dataout_7_), .C(mac1_reset_bF_buf0), .Y(_787_) );
NAND3X1 NAND3X1_246 ( .A(_780_), .B(_784_), .C(_787_), .Y(_789_) );
AOI21X1 AOI21X1_44 ( .A(_776_), .B(_778_), .C(_713_), .Y(_790_) );
AOI21X1 AOI21X1_45 ( .A(_769_), .B(_772_), .C(_712_), .Y(_791_) );
AND2X2 AND2X2_40 ( .A(_783_), .B(_781_), .Y(_792_) );
OAI21X1 OAI21X1_84 ( .A(_781_), .B(_783_), .C(_745_), .Y(_793_) );
OAI22X1 OAI22X1_52 ( .A(_790_), .B(_791_), .C(_793_), .D(_792_), .Y(_794_) );
NAND2X1 NAND2X1_115 ( .A(_794_), .B(_789_), .Y(_487__7_) );
DFFPOSX1 DFFPOSX1_14 ( .CLK(clk_bF_buf0), .D(_487__0_), .Q(mac1_dataout_0_) );
DFFPOSX1 DFFPOSX1_15 ( .CLK(clk_bF_buf6), .D(_487__1_), .Q(mac1_dataout_1_) );
DFFPOSX1 DFFPOSX1_16 ( .CLK(clk_bF_buf5), .D(_487__2_), .Q(mac1_dataout_2_) );
DFFPOSX1 DFFPOSX1_17 ( .CLK(clk_bF_buf4), .D(_487__3_), .Q(mac1_dataout_3_) );
DFFPOSX1 DFFPOSX1_18 ( .CLK(clk_bF_buf3), .D(_487__4_), .Q(mac1_dataout_4_) );
DFFPOSX1 DFFPOSX1_19 ( .CLK(clk_bF_buf2), .D(_487__5_), .Q(mac1_dataout_5_) );
DFFPOSX1 DFFPOSX1_20 ( .CLK(clk_bF_buf1), .D(_487__6_), .Q(mac1_dataout_6_) );
DFFPOSX1 DFFPOSX1_21 ( .CLK(clk_bF_buf0), .D(_487__7_), .Q(mac1_dataout_7_) );
INVX1 INVX1_181 ( .A(reg1_dataout_0_), .Y(_855_) );
NAND2X1 NAND2X1_116 ( .A(din[0]), .B(vdd), .Y(_856_) );
OAI21X1 OAI21X1_85 ( .A(vdd), .B(_855_), .C(_856_), .Y(_853__0_) );
INVX1 INVX1_182 ( .A(reg1_dataout_1_), .Y(_857_) );
NAND2X1 NAND2X1_117 ( .A(vdd), .B(din[1]), .Y(_858_) );
OAI21X1 OAI21X1_86 ( .A(vdd), .B(_857_), .C(_858_), .Y(_853__1_) );
INVX1 INVX1_183 ( .A(reg1_dataout_2_), .Y(_859_) );
NAND2X1 NAND2X1_118 ( .A(vdd), .B(din[2]), .Y(_860_) );
OAI21X1 OAI21X1_87 ( .A(vdd), .B(_859_), .C(_860_), .Y(_853__2_) );
INVX1 INVX1_184 ( .A(reg1_dataout_3_), .Y(_861_) );
NAND2X1 NAND2X1_119 ( .A(vdd), .B(din[3]), .Y(_862_) );
OAI21X1 OAI21X1_88 ( .A(vdd), .B(_861_), .C(_862_), .Y(_853__3_) );
INVX1 INVX1_185 ( .A(reg1_dataout_4_), .Y(_863_) );
NAND2X1 NAND2X1_120 ( .A(vdd), .B(din[4]), .Y(_864_) );
OAI21X1 OAI21X1_89 ( .A(vdd), .B(_863_), .C(_864_), .Y(_853__4_) );
INVX1 INVX1_186 ( .A(reg1_dataout_5_), .Y(_865_) );
NAND2X1 NAND2X1_121 ( .A(vdd), .B(din[5]), .Y(_866_) );
OAI21X1 OAI21X1_90 ( .A(vdd), .B(_865_), .C(_866_), .Y(_853__5_) );
INVX1 INVX1_187 ( .A(reg1_dataout_6_), .Y(_867_) );
NAND2X1 NAND2X1_122 ( .A(vdd), .B(din[6]), .Y(_868_) );
OAI21X1 OAI21X1_91 ( .A(vdd), .B(_867_), .C(_868_), .Y(_853__6_) );
INVX1 INVX1_188 ( .A(reg1_dataout_7_), .Y(_869_) );
NAND2X1 NAND2X1_123 ( .A(vdd), .B(din[7]), .Y(_870_) );
OAI21X1 OAI21X1_92 ( .A(vdd), .B(_869_), .C(_870_), .Y(_853__7_) );
INVX1 INVX1_189 ( .A(rst_bF_buf5), .Y(_854_) );
DFFSR DFFSR_257 ( .CLK(clk2_clkout_bF_buf35), .D(_853__0_), .Q(reg1_dataout_0_), .R(_854_), .S(vdd) );
DFFSR DFFSR_258 ( .CLK(clk2_clkout_bF_buf34), .D(_853__1_), .Q(reg1_dataout_1_), .R(_854_), .S(vdd) );
DFFSR DFFSR_259 ( .CLK(clk2_clkout_bF_buf33), .D(_853__2_), .Q(reg1_dataout_2_), .R(_854_), .S(vdd) );
DFFSR DFFSR_260 ( .CLK(clk2_clkout_bF_buf32), .D(_853__3_), .Q(reg1_dataout_3_), .R(_854_), .S(vdd) );
DFFSR DFFSR_261 ( .CLK(clk2_clkout_bF_buf31), .D(_853__4_), .Q(reg1_dataout_4_), .R(_854_), .S(vdd) );
DFFSR DFFSR_262 ( .CLK(clk2_clkout_bF_buf30), .D(_853__5_), .Q(reg1_dataout_5_), .R(_854_), .S(vdd) );
DFFSR DFFSR_263 ( .CLK(clk2_clkout_bF_buf29), .D(_853__6_), .Q(reg1_dataout_6_), .R(_854_), .S(vdd) );
DFFSR DFFSR_264 ( .CLK(clk2_clkout_bF_buf28), .D(_853__7_), .Q(reg1_dataout_7_), .R(_854_), .S(vdd) );
INVX1 INVX1_190 ( .A(reg2_dataout_0_), .Y(_873_) );
NAND2X1 NAND2X1_124 ( .A(mac1_dataout_0_), .B(mac1_reset_bF_buf3), .Y(_874_) );
OAI21X1 OAI21X1_93 ( .A(mac1_reset_bF_buf2), .B(_873_), .C(_874_), .Y(_871__0_) );
INVX1 INVX1_191 ( .A(reg2_dataout_1_), .Y(_875_) );
NAND2X1 NAND2X1_125 ( .A(mac1_reset_bF_buf1), .B(mac1_dataout_1_), .Y(_876_) );
OAI21X1 OAI21X1_94 ( .A(mac1_reset_bF_buf0), .B(_875_), .C(_876_), .Y(_871__1_) );
INVX1 INVX1_192 ( .A(reg2_dataout_2_), .Y(_877_) );
NAND2X1 NAND2X1_126 ( .A(mac1_reset_bF_buf3), .B(mac1_dataout_2_), .Y(_878_) );
OAI21X1 OAI21X1_95 ( .A(mac1_reset_bF_buf2), .B(_877_), .C(_878_), .Y(_871__2_) );
INVX1 INVX1_193 ( .A(reg2_dataout_3_), .Y(_879_) );
NAND2X1 NAND2X1_127 ( .A(mac1_reset_bF_buf1), .B(mac1_dataout_3_), .Y(_880_) );
OAI21X1 OAI21X1_96 ( .A(mac1_reset_bF_buf0), .B(_879_), .C(_880_), .Y(_871__3_) );
INVX1 INVX1_194 ( .A(reg2_dataout_4_), .Y(_881_) );
NAND2X1 NAND2X1_128 ( .A(mac1_reset_bF_buf3), .B(mac1_dataout_4_), .Y(_882_) );
OAI21X1 OAI21X1_97 ( .A(mac1_reset_bF_buf2), .B(_881_), .C(_882_), .Y(_871__4_) );
INVX1 INVX1_195 ( .A(reg2_dataout_5_), .Y(_883_) );
NAND2X1 NAND2X1_129 ( .A(mac1_reset_bF_buf1), .B(mac1_dataout_5_), .Y(_884_) );
OAI21X1 OAI21X1_98 ( .A(mac1_reset_bF_buf0), .B(_883_), .C(_884_), .Y(_871__5_) );
INVX1 INVX1_196 ( .A(reg2_dataout_6_), .Y(_885_) );
NAND2X1 NAND2X1_130 ( .A(mac1_reset_bF_buf3), .B(mac1_dataout_6_), .Y(_886_) );
OAI21X1 OAI21X1_99 ( .A(mac1_reset_bF_buf2), .B(_885_), .C(_886_), .Y(_871__6_) );
INVX1 INVX1_197 ( .A(reg2_dataout_7_), .Y(_887_) );
NAND2X1 NAND2X1_131 ( .A(mac1_reset_bF_buf1), .B(mac1_dataout_7_), .Y(_888_) );
OAI21X1 OAI21X1_100 ( .A(mac1_reset_bF_buf0), .B(_887_), .C(_888_), .Y(_871__7_) );
INVX1 INVX1_198 ( .A(rst_bF_buf4), .Y(_872_) );
DFFSR DFFSR_265 ( .CLK(clk_bF_buf6), .D(_871__0_), .Q(reg2_dataout_0_), .R(_872_), .S(vdd) );
DFFSR DFFSR_266 ( .CLK(clk_bF_buf5), .D(_871__1_), .Q(reg2_dataout_1_), .R(_872_), .S(vdd) );
DFFSR DFFSR_267 ( .CLK(clk_bF_buf4), .D(_871__2_), .Q(reg2_dataout_2_), .R(_872_), .S(vdd) );
DFFSR DFFSR_268 ( .CLK(clk_bF_buf3), .D(_871__3_), .Q(reg2_dataout_3_), .R(_872_), .S(vdd) );
DFFSR DFFSR_269 ( .CLK(clk_bF_buf2), .D(_871__4_), .Q(reg2_dataout_4_), .R(_872_), .S(vdd) );
DFFSR DFFSR_270 ( .CLK(clk_bF_buf1), .D(_871__5_), .Q(reg2_dataout_5_), .R(_872_), .S(vdd) );
DFFSR DFFSR_271 ( .CLK(clk_bF_buf0), .D(_871__6_), .Q(reg2_dataout_6_), .R(_872_), .S(vdd) );
DFFSR DFFSR_272 ( .CLK(clk_bF_buf6), .D(_871__7_), .Q(reg2_dataout_7_), .R(_872_), .S(vdd) );
INVX1 INVX1_199 ( .A(reg3_dataout_0_), .Y(_891_) );
NAND2X1 NAND2X1_132 ( .A(reg2_dataout_0_), .B(vdd), .Y(_892_) );
OAI21X1 OAI21X1_101 ( .A(vdd), .B(_891_), .C(_892_), .Y(_889__0_) );
INVX1 INVX1_200 ( .A(reg3_dataout_1_), .Y(_893_) );
NAND2X1 NAND2X1_133 ( .A(vdd), .B(reg2_dataout_1_), .Y(_894_) );
OAI21X1 OAI21X1_102 ( .A(vdd), .B(_893_), .C(_894_), .Y(_889__1_) );
INVX1 INVX1_201 ( .A(reg3_dataout_2_), .Y(_895_) );
NAND2X1 NAND2X1_134 ( .A(vdd), .B(reg2_dataout_2_), .Y(_896_) );
OAI21X1 OAI21X1_103 ( .A(vdd), .B(_895_), .C(_896_), .Y(_889__2_) );
INVX1 INVX1_202 ( .A(reg3_dataout_3_), .Y(_897_) );
NAND2X1 NAND2X1_135 ( .A(vdd), .B(reg2_dataout_3_), .Y(_898_) );
OAI21X1 OAI21X1_104 ( .A(vdd), .B(_897_), .C(_898_), .Y(_889__3_) );
INVX1 INVX1_203 ( .A(reg3_dataout_4_), .Y(_899_) );
NAND2X1 NAND2X1_136 ( .A(vdd), .B(reg2_dataout_4_), .Y(_900_) );
OAI21X1 OAI21X1_105 ( .A(vdd), .B(_899_), .C(_900_), .Y(_889__4_) );
INVX1 INVX1_204 ( .A(reg3_dataout_5_), .Y(_901_) );
NAND2X1 NAND2X1_137 ( .A(vdd), .B(reg2_dataout_5_), .Y(_902_) );
OAI21X1 OAI21X1_106 ( .A(vdd), .B(_901_), .C(_902_), .Y(_889__5_) );
INVX1 INVX1_205 ( .A(reg3_dataout_6_), .Y(_903_) );
NAND2X1 NAND2X1_138 ( .A(vdd), .B(reg2_dataout_6_), .Y(_904_) );
OAI21X1 OAI21X1_107 ( .A(vdd), .B(_903_), .C(_904_), .Y(_889__6_) );
INVX1 INVX1_206 ( .A(reg3_dataout_7_), .Y(_905_) );
NAND2X1 NAND2X1_139 ( .A(vdd), .B(reg2_dataout_7_), .Y(_906_) );
OAI21X1 OAI21X1_108 ( .A(vdd), .B(_905_), .C(_906_), .Y(_889__7_) );
INVX1 INVX1_207 ( .A(rst_bF_buf3), .Y(_890_) );
DFFSR DFFSR_273 ( .CLK(clk2_clkout_bF_buf27), .D(_889__0_), .Q(reg3_dataout_0_), .R(_890_), .S(vdd) );
DFFSR DFFSR_274 ( .CLK(clk2_clkout_bF_buf26), .D(_889__1_), .Q(reg3_dataout_1_), .R(_890_), .S(vdd) );
DFFSR DFFSR_275 ( .CLK(clk2_clkout_bF_buf25), .D(_889__2_), .Q(reg3_dataout_2_), .R(_890_), .S(vdd) );
DFFSR DFFSR_276 ( .CLK(clk2_clkout_bF_buf24), .D(_889__3_), .Q(reg3_dataout_3_), .R(_890_), .S(vdd) );
DFFSR DFFSR_277 ( .CLK(clk2_clkout_bF_buf23), .D(_889__4_), .Q(reg3_dataout_4_), .R(_890_), .S(vdd) );
DFFSR DFFSR_278 ( .CLK(clk2_clkout_bF_buf22), .D(_889__5_), .Q(reg3_dataout_5_), .R(_890_), .S(vdd) );
DFFSR DFFSR_279 ( .CLK(clk2_clkout_bF_buf21), .D(_889__6_), .Q(reg3_dataout_6_), .R(_890_), .S(vdd) );
DFFSR DFFSR_280 ( .CLK(clk2_clkout_bF_buf20), .D(_889__7_), .Q(reg3_dataout_7_), .R(_890_), .S(vdd) );
INVX1 INVX1_208 ( .A(vdd), .Y(_923_) );
NAND2X1 NAND2X1_140 ( .A(ret2_rf_13_), .B(_923_), .Y(_924_) );
NAND2X1 NAND2X1_141 ( .A(ret2_rf_12_), .B(vdd), .Y(_925_) );
AOI21X1 AOI21X1_46 ( .A(_924_), .B(_925_), .C(rst_bF_buf2), .Y(_912_) );
NAND2X1 NAND2X1_142 ( .A(ret2_rf_14_), .B(_923_), .Y(_926_) );
NAND2X1 NAND2X1_143 ( .A(ret2_rf_13_), .B(vdd), .Y(_927_) );
AOI21X1 AOI21X1_47 ( .A(_926_), .B(_927_), .C(rst_bF_buf1), .Y(_913_) );
NAND2X1 NAND2X1_144 ( .A(ret2_rf_12_), .B(_923_), .Y(_928_) );
NAND2X1 NAND2X1_145 ( .A(vdd), .B(ret2_rf_11_), .Y(_929_) );
AOI21X1 AOI21X1_48 ( .A(_928_), .B(_929_), .C(rst_bF_buf0), .Y(_911_) );
NAND2X1 NAND2X1_146 ( .A(ret2_rf_11_), .B(_923_), .Y(_930_) );
NAND2X1 NAND2X1_147 ( .A(vdd), .B(ret2_rf_10_), .Y(_931_) );
AOI21X1 AOI21X1_49 ( .A(_930_), .B(_931_), .C(rst_bF_buf5), .Y(_910_) );
NAND2X1 NAND2X1_148 ( .A(ret2_rf_10_), .B(_923_), .Y(_932_) );
NAND2X1 NAND2X1_149 ( .A(vdd), .B(ret2_rf_9_), .Y(_933_) );
AOI21X1 AOI21X1_50 ( .A(_932_), .B(_933_), .C(rst_bF_buf4), .Y(_909_) );
NAND2X1 NAND2X1_150 ( .A(ret2_rf_9_), .B(_923_), .Y(_934_) );
NAND2X1 NAND2X1_151 ( .A(vdd), .B(ret2_rf_8_), .Y(_935_) );
AOI21X1 AOI21X1_51 ( .A(_934_), .B(_935_), .C(rst_bF_buf3), .Y(_922_) );
NAND2X1 NAND2X1_152 ( .A(ret2_rf_8_), .B(_923_), .Y(_936_) );
NAND2X1 NAND2X1_153 ( .A(vdd), .B(ret2_rf_7_), .Y(_937_) );
AOI21X1 AOI21X1_52 ( .A(_936_), .B(_937_), .C(rst_bF_buf2), .Y(_921_) );
NAND2X1 NAND2X1_154 ( .A(ret2_rf_7_), .B(_923_), .Y(_938_) );
NAND2X1 NAND2X1_155 ( .A(vdd), .B(ret2_rf_6_), .Y(_939_) );
AOI21X1 AOI21X1_53 ( .A(_938_), .B(_939_), .C(rst_bF_buf1), .Y(_920_) );
NAND2X1 NAND2X1_156 ( .A(ret2_rf_6_), .B(_923_), .Y(_940_) );
NAND2X1 NAND2X1_157 ( .A(vdd), .B(ret2_rf_5_), .Y(_941_) );
AOI21X1 AOI21X1_54 ( .A(_940_), .B(_941_), .C(rst_bF_buf0), .Y(_919_) );
NAND2X1 NAND2X1_158 ( .A(ret2_rf_5_), .B(_923_), .Y(_942_) );
NAND2X1 NAND2X1_159 ( .A(vdd), .B(ret2_rf_4_), .Y(_943_) );
AOI21X1 AOI21X1_55 ( .A(_942_), .B(_943_), .C(rst_bF_buf5), .Y(_918_) );
NAND2X1 NAND2X1_160 ( .A(ret2_rf_4_), .B(_923_), .Y(_944_) );
NAND2X1 NAND2X1_161 ( .A(vdd), .B(ret2_rf_3_), .Y(_945_) );
AOI21X1 AOI21X1_56 ( .A(_944_), .B(_945_), .C(rst_bF_buf4), .Y(_917_) );
NAND2X1 NAND2X1_162 ( .A(ret2_rf_3_), .B(_923_), .Y(_946_) );
NAND2X1 NAND2X1_163 ( .A(vdd), .B(ret2_rf_2_), .Y(_947_) );
AOI21X1 AOI21X1_57 ( .A(_946_), .B(_947_), .C(rst_bF_buf3), .Y(_916_) );
NAND2X1 NAND2X1_164 ( .A(ret2_rf_2_), .B(_923_), .Y(_948_) );
NAND2X1 NAND2X1_165 ( .A(vdd), .B(ret2_rf_1_), .Y(_949_) );
AOI21X1 AOI21X1_58 ( .A(_948_), .B(_949_), .C(rst_bF_buf2), .Y(_915_) );
NAND2X1 NAND2X1_166 ( .A(ret2_rf_1_), .B(_923_), .Y(_950_) );
NAND2X1 NAND2X1_167 ( .A(vdd), .B(ret2_rf_0_), .Y(_951_) );
AOI21X1 AOI21X1_59 ( .A(_950_), .B(_951_), .C(rst_bF_buf1), .Y(_914_) );
NAND2X1 NAND2X1_168 ( .A(ret2_rf_0_), .B(_923_), .Y(_952_) );
NAND2X1 NAND2X1_169 ( .A(vdd), .B(comp_dataout), .Y(_953_) );
AOI21X1 AOI21X1_60 ( .A(_952_), .B(_953_), .C(rst_bF_buf0), .Y(_908_) );
NAND2X1 NAND2X1_170 ( .A(vdd), .B(ret2_rf_14_), .Y(_954_) );
NOR2X1 NOR2X1_74 ( .A(rst_bF_buf5), .B(_954_), .Y(_907_) );
DFFPOSX1 DFFPOSX1_22 ( .CLK(clk_bF_buf5), .D(_907_), .Q(mac1_reset) );
DFFPOSX1 DFFPOSX1_23 ( .CLK(clk_bF_buf4), .D(_917_), .Q(ret2_rf_4_) );
DFFPOSX1 DFFPOSX1_24 ( .CLK(clk_bF_buf3), .D(_914_), .Q(ret2_rf_1_) );
DFFPOSX1 DFFPOSX1_25 ( .CLK(clk_bF_buf2), .D(_908_), .Q(ret2_rf_0_) );
DFFPOSX1 DFFPOSX1_26 ( .CLK(clk_bF_buf1), .D(_919_), .Q(ret2_rf_6_) );
DFFPOSX1 DFFPOSX1_27 ( .CLK(clk_bF_buf0), .D(_922_), .Q(ret2_rf_9_) );
DFFPOSX1 DFFPOSX1_28 ( .CLK(clk_bF_buf6), .D(_909_), .Q(ret2_rf_10_) );
DFFPOSX1 DFFPOSX1_29 ( .CLK(clk_bF_buf5), .D(_916_), .Q(ret2_rf_3_) );
DFFPOSX1 DFFPOSX1_30 ( .CLK(clk_bF_buf4), .D(_920_), .Q(ret2_rf_7_) );
DFFPOSX1 DFFPOSX1_31 ( .CLK(clk_bF_buf3), .D(_921_), .Q(ret2_rf_8_) );
DFFPOSX1 DFFPOSX1_32 ( .CLK(clk_bF_buf2), .D(_915_), .Q(ret2_rf_2_) );
DFFPOSX1 DFFPOSX1_33 ( .CLK(clk_bF_buf1), .D(_918_), .Q(ret2_rf_5_) );
DFFPOSX1 DFFPOSX1_34 ( .CLK(clk_bF_buf0), .D(_910_), .Q(ret2_rf_11_) );
DFFPOSX1 DFFPOSX1_35 ( .CLK(clk_bF_buf6), .D(_911_), .Q(ret2_rf_12_) );
DFFPOSX1 DFFPOSX1_36 ( .CLK(clk_bF_buf5), .D(_912_), .Q(ret2_rf_13_) );
DFFPOSX1 DFFPOSX1_37 ( .CLK(clk_bF_buf4), .D(_913_), .Q(ret2_rf_14_) );
NOR2X1 NOR2X1_75 ( .A(counterup_counter_0_bF_buf2_), .B(rst_bF_buf4), .Y(_955__0_) );
INVX1 INVX1_209 ( .A(rst_bF_buf3), .Y(_956_) );
OAI21X1 OAI21X1_109 ( .A(counterup_counter_0_bF_buf1_), .B(counterup_counter_1_), .C(_956_), .Y(_957_) );
AOI21X1 AOI21X1_61 ( .A(counterup_counter_0_bF_buf0_), .B(counterup_counter_1_), .C(_957_), .Y(_955__1_) );
AOI21X1 AOI21X1_62 ( .A(counterup_counter_0_bF_buf3_), .B(counterup_counter_1_), .C(counterup_counter_2_), .Y(_958_) );
NAND3X1 NAND3X1_247 ( .A(counterup_counter_0_bF_buf2_), .B(counterup_counter_1_), .C(counterup_counter_2_), .Y(_959_) );
NAND2X1 NAND2X1_171 ( .A(_956_), .B(_959_), .Y(_960_) );
NOR2X1 NOR2X1_76 ( .A(_958_), .B(_960_), .Y(_955__2_) );
INVX1 INVX1_210 ( .A(counterup_counter_3_), .Y(_961_) );
OAI21X1 OAI21X1_110 ( .A(_961_), .B(_959_), .C(_956_), .Y(_962_) );
AOI21X1 AOI21X1_63 ( .A(_961_), .B(_959_), .C(_962_), .Y(_955__3_) );
NOR3X1 NOR3X1_6 ( .A(rst_bF_buf2), .B(_961_), .C(_959_), .Y(_955__4_) );
DFFPOSX1 DFFPOSX1_38 ( .CLK(clk_bF_buf3), .D(_955__0_), .Q(rom1_data_0_) );
DFFPOSX1 DFFPOSX1_39 ( .CLK(clk_bF_buf2), .D(_955__1_), .Q(rom1_data_1_) );
DFFPOSX1 DFFPOSX1_40 ( .CLK(clk_bF_buf1), .D(_955__2_), .Q(rom1_data_2_) );
DFFPOSX1 DFFPOSX1_41 ( .CLK(clk_bF_buf0), .D(_955__3_), .Q(rom1_data_3_) );
DFFPOSX1 DFFPOSX1_42 ( .CLK(clk_bF_buf6), .D(_955__4_), .Q(rom1_data_4_) );
NAND2X1 NAND2X1_172 ( .A(asr1_dataout_0_), .B(asr2_dataout_0_), .Y(_964_) );
INVX1 INVX1_211 ( .A(_964_), .Y(_965_) );
INVX1 INVX1_212 ( .A(rst_bF_buf1), .Y(_966_) );
OAI21X1 OAI21X1_111 ( .A(asr1_dataout_0_), .B(asr2_dataout_0_), .C(_966_), .Y(_967_) );
NOR2X1 NOR2X1_77 ( .A(_965_), .B(_967_), .Y(_963__0_) );
XOR2X1 XOR2X1_9 ( .A(asr1_dataout_1_), .B(asr2_dataout_1_), .Y(_968_) );
AND2X2 AND2X2_41 ( .A(_968_), .B(_965_), .Y(_969_) );
OAI21X1 OAI21X1_112 ( .A(_965_), .B(_968_), .C(_966_), .Y(_970_) );
OR2X2 OR2X2_5 ( .A(_969_), .B(_970_), .Y(_971_) );
INVX1 INVX1_213 ( .A(_971_), .Y(_963__1_) );
NOR2X1 NOR2X1_78 ( .A(asr1_dataout_1_), .B(asr2_dataout_1_), .Y(_972_) );
NAND2X1 NAND2X1_173 ( .A(asr1_dataout_1_), .B(asr2_dataout_1_), .Y(_973_) );
OAI21X1 OAI21X1_113 ( .A(_964_), .B(_972_), .C(_973_), .Y(_974_) );
XOR2X1 XOR2X1_10 ( .A(asr1_dataout_2_), .B(asr2_dataout_2_), .Y(_975_) );
OAI21X1 OAI21X1_114 ( .A(_975_), .B(_974_), .C(_966_), .Y(_976_) );
AOI21X1 AOI21X1_64 ( .A(_974_), .B(_975_), .C(_976_), .Y(_963__2_) );
XOR2X1 XOR2X1_11 ( .A(asr1_dataout_3_), .B(asr2_dataout_3_), .Y(_977_) );
AND2X2 AND2X2_42 ( .A(asr1_dataout_2_), .B(asr2_dataout_2_), .Y(_978_) );
AOI21X1 AOI21X1_65 ( .A(_974_), .B(_975_), .C(_978_), .Y(_979_) );
XOR2X1 XOR2X1_12 ( .A(_979_), .B(_977_), .Y(_980_) );
NOR2X1 NOR2X1_79 ( .A(rst_bF_buf0), .B(_980_), .Y(_963__3_) );
NAND3X1 NAND3X1_248 ( .A(_975_), .B(_977_), .C(_974_), .Y(_981_) );
INVX1 INVX1_214 ( .A(asr1_dataout_3_), .Y(_982_) );
INVX1 INVX1_215 ( .A(asr2_dataout_3_), .Y(_983_) );
NAND2X1 NAND2X1_174 ( .A(_982_), .B(_983_), .Y(_984_) );
NOR2X1 NOR2X1_80 ( .A(_982_), .B(_983_), .Y(_985_) );
AOI21X1 AOI21X1_66 ( .A(_978_), .B(_984_), .C(_985_), .Y(_986_) );
NAND2X1 NAND2X1_175 ( .A(_986_), .B(_981_), .Y(_987_) );
XOR2X1 XOR2X1_13 ( .A(asr1_dataout_4_), .B(asr2_dataout_4_), .Y(_988_) );
OAI21X1 OAI21X1_115 ( .A(_988_), .B(_987_), .C(_966_), .Y(_989_) );
AOI21X1 AOI21X1_67 ( .A(_987_), .B(_988_), .C(_989_), .Y(_963__4_) );
XOR2X1 XOR2X1_14 ( .A(asr1_dataout_5_), .B(asr2_dataout_5_), .Y(_990_) );
NAND2X1 NAND2X1_176 ( .A(_988_), .B(_990_), .Y(_991_) );
AOI21X1 AOI21X1_68 ( .A(_981_), .B(_986_), .C(_991_), .Y(_992_) );
INVX1 INVX1_216 ( .A(asr1_dataout_4_), .Y(_993_) );
INVX1 INVX1_217 ( .A(asr2_dataout_4_), .Y(_994_) );
NAND2X1 NAND2X1_177 ( .A(_988_), .B(_987_), .Y(_995_) );
OAI21X1 OAI21X1_116 ( .A(_993_), .B(_994_), .C(_995_), .Y(_996_) );
NOR2X1 NOR2X1_81 ( .A(_993_), .B(_994_), .Y(_997_) );
AOI21X1 AOI21X1_69 ( .A(_990_), .B(_997_), .C(rst_bF_buf5), .Y(_998_) );
OAI21X1 OAI21X1_117 ( .A(_990_), .B(_996_), .C(_998_), .Y(_999_) );
NOR2X1 NOR2X1_82 ( .A(_992_), .B(_999_), .Y(_963__5_) );
NAND2X1 NAND2X1_178 ( .A(asr1_dataout_5_), .B(asr2_dataout_5_), .Y(_1000_) );
NAND2X1 NAND2X1_179 ( .A(_997_), .B(_990_), .Y(_1001_) );
NAND2X1 NAND2X1_180 ( .A(_1000_), .B(_1001_), .Y(_1002_) );
OR2X2 OR2X2_6 ( .A(_992_), .B(_1002_), .Y(_1003_) );
XOR2X1 XOR2X1_15 ( .A(asr1_dataout_6_), .B(asr2_dataout_6_), .Y(_1004_) );
OAI21X1 OAI21X1_118 ( .A(_1004_), .B(_1003_), .C(_966_), .Y(_1005_) );
AOI21X1 AOI21X1_70 ( .A(_1003_), .B(_1004_), .C(_1005_), .Y(_963__6_) );
NAND2X1 NAND2X1_181 ( .A(asr1_dataout_6_), .B(asr2_dataout_6_), .Y(_1006_) );
OAI21X1 OAI21X1_119 ( .A(_1002_), .B(_992_), .C(_1004_), .Y(_1007_) );
XNOR2X1 XNOR2X1_4 ( .A(asr1_dataout_7_), .B(asr2_dataout_7_), .Y(_1008_) );
AOI21X1 AOI21X1_71 ( .A(_1007_), .B(_1006_), .C(_1008_), .Y(_1009_) );
NAND3X1 NAND3X1_249 ( .A(_1006_), .B(_1008_), .C(_1007_), .Y(_1010_) );
NAND2X1 NAND2X1_182 ( .A(_966_), .B(_1010_), .Y(_1011_) );
NOR2X1 NOR2X1_83 ( .A(_1009_), .B(_1011_), .Y(_963__7_) );
DFFPOSX1 DFFPOSX1_43 ( .CLK(clk_bF_buf5), .D(_963__0_), .Q(sumador_res_0_) );
DFFPOSX1 DFFPOSX1_44 ( .CLK(clk_bF_buf4), .D(_963__1_), .Q(sumador_res_1_) );
DFFPOSX1 DFFPOSX1_45 ( .CLK(clk_bF_buf3), .D(_963__2_), .Q(sumador_res_2_) );
DFFPOSX1 DFFPOSX1_46 ( .CLK(clk_bF_buf2), .D(_963__3_), .Q(sumador_res_3_) );
DFFPOSX1 DFFPOSX1_47 ( .CLK(clk_bF_buf1), .D(_963__4_), .Q(sumador_res_4_) );
DFFPOSX1 DFFPOSX1_48 ( .CLK(clk_bF_buf0), .D(_963__5_), .Q(sumador_res_5_) );
DFFPOSX1 DFFPOSX1_49 ( .CLK(clk_bF_buf6), .D(_963__6_), .Q(sumador_res_6_) );
DFFPOSX1 DFFPOSX1_50 ( .CLK(clk_bF_buf5), .D(_963__7_), .Q(sumador_res_7_) );
BUFX2 BUFX2_79 ( .A(gnd), .Y(_955__5_) );
BUFX2 BUFX2_80 ( .A(gnd), .Y(_955__6_) );
BUFX2 BUFX2_81 ( .A(gnd), .Y(_955__7_) );
BUFX2 BUFX2_82 ( .A(asr1_en_0_), .Y(asr1_rom_15__0_) );
BUFX2 BUFX2_83 ( .A(asr1_en_1_), .Y(asr1_rom_15__1_) );
BUFX2 BUFX2_84 ( .A(asr1_en_2_), .Y(asr1_rom_15__2_) );
BUFX2 BUFX2_85 ( .A(asr1_en_3_), .Y(asr1_rom_15__3_) );
BUFX2 BUFX2_86 ( .A(asr1_en_4_), .Y(asr1_rom_15__4_) );
BUFX2 BUFX2_87 ( .A(asr1_en_5_), .Y(asr1_rom_15__5_) );
BUFX2 BUFX2_88 ( .A(asr1_en_6_), .Y(asr1_rom_15__6_) );
BUFX2 BUFX2_89 ( .A(asr1_en_7_), .Y(asr1_rom_15__7_) );
BUFX2 BUFX2_90 ( .A(asr2_en_0_), .Y(asr2_rom_15__0_) );
BUFX2 BUFX2_91 ( .A(asr2_en_1_), .Y(asr2_rom_15__1_) );
BUFX2 BUFX2_92 ( .A(asr2_en_2_), .Y(asr2_rom_15__2_) );
BUFX2 BUFX2_93 ( .A(asr2_en_3_), .Y(asr2_rom_15__3_) );
BUFX2 BUFX2_94 ( .A(asr2_en_4_), .Y(asr2_rom_15__4_) );
BUFX2 BUFX2_95 ( .A(asr2_en_5_), .Y(asr2_rom_15__5_) );
BUFX2 BUFX2_96 ( .A(asr2_en_6_), .Y(asr2_rom_15__6_) );
BUFX2 BUFX2_97 ( .A(asr2_en_7_), .Y(asr2_rom_15__7_) );
BUFX2 BUFX2_98 ( .A(gnd), .Y(rom1_data_5_) );
BUFX2 BUFX2_99 ( .A(gnd), .Y(rom1_data_6_) );
BUFX2 BUFX2_100 ( .A(gnd), .Y(rom1_data_7_) );
endmodule
